magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 86 368 116 536
rect 193 368 223 592
rect 283 368 313 592
rect 428 368 458 568
rect 512 368 542 568
rect 620 368 650 568
<< nmoslvt >>
rect 98 112 128 222
rect 200 74 230 222
rect 286 74 316 222
rect 431 94 461 222
rect 531 94 561 222
rect 645 94 675 222
<< ndiff >>
rect 41 184 98 222
rect 41 150 53 184
rect 87 150 98 184
rect 41 112 98 150
rect 128 131 200 222
rect 128 112 155 131
rect 143 97 155 112
rect 189 97 200 131
rect 143 74 200 97
rect 230 210 286 222
rect 230 176 241 210
rect 275 176 286 210
rect 230 120 286 176
rect 230 86 241 120
rect 275 86 286 120
rect 230 74 286 86
rect 316 147 431 222
rect 316 113 363 147
rect 397 113 431 147
rect 316 94 431 113
rect 461 210 531 222
rect 461 176 486 210
rect 520 176 531 210
rect 461 140 531 176
rect 461 106 486 140
rect 520 106 531 140
rect 461 94 531 106
rect 561 146 645 222
rect 561 112 586 146
rect 620 112 645 146
rect 561 94 645 112
rect 675 210 732 222
rect 675 176 686 210
rect 720 176 732 210
rect 675 140 732 176
rect 675 106 686 140
rect 720 106 732 140
rect 675 94 732 106
rect 316 74 366 94
<< pdiff >>
rect 331 592 410 594
rect 134 573 193 592
rect 134 539 146 573
rect 180 539 193 573
rect 134 536 193 539
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 440 86 490
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 368 193 536
rect 223 414 283 592
rect 223 380 236 414
rect 270 380 283 414
rect 223 368 283 380
rect 313 582 410 592
rect 313 548 353 582
rect 387 568 410 582
rect 387 548 428 568
rect 313 368 428 548
rect 458 368 512 568
rect 542 368 620 568
rect 650 560 709 568
rect 650 526 663 560
rect 697 526 709 560
rect 650 492 709 526
rect 650 458 663 492
rect 697 458 709 492
rect 650 368 709 458
<< ndiffc >>
rect 53 150 87 184
rect 155 97 189 131
rect 241 176 275 210
rect 241 86 275 120
rect 363 113 397 147
rect 486 176 520 210
rect 486 106 520 140
rect 586 112 620 146
rect 686 176 720 210
rect 686 106 720 140
<< pdiffc >>
rect 146 539 180 573
rect 39 490 73 524
rect 39 406 73 440
rect 236 380 270 414
rect 353 548 387 582
rect 663 526 697 560
rect 663 458 697 492
<< poly >>
rect 193 592 223 618
rect 283 592 313 618
rect 86 536 116 562
rect 428 568 458 594
rect 512 568 542 594
rect 620 568 650 594
rect 86 353 116 368
rect 193 353 223 368
rect 283 353 313 368
rect 428 353 458 368
rect 512 353 542 368
rect 620 353 650 368
rect 83 338 116 353
rect 83 326 113 338
rect 21 310 113 326
rect 21 276 37 310
rect 71 290 113 310
rect 190 290 226 353
rect 280 326 316 353
rect 425 336 461 353
rect 509 336 545 353
rect 617 345 653 353
rect 280 310 347 326
rect 280 290 297 310
rect 71 276 128 290
rect 21 260 128 276
rect 190 276 297 290
rect 331 276 347 310
rect 190 260 347 276
rect 395 320 461 336
rect 395 286 411 320
rect 445 286 461 320
rect 395 270 461 286
rect 503 320 569 336
rect 503 286 519 320
rect 553 286 569 320
rect 503 270 569 286
rect 617 320 683 345
rect 617 286 633 320
rect 667 286 683 320
rect 617 270 683 286
rect 98 222 128 260
rect 200 222 230 260
rect 286 222 316 260
rect 431 222 461 270
rect 531 222 561 270
rect 645 222 675 270
rect 98 86 128 112
rect 200 48 230 74
rect 286 48 316 74
rect 431 68 461 94
rect 531 68 561 94
rect 645 68 675 94
<< polycont >>
rect 37 276 71 310
rect 297 276 331 310
rect 411 286 445 320
rect 519 286 553 320
rect 633 286 667 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 130 573 196 649
rect 23 524 89 540
rect 130 539 146 573
rect 180 539 196 573
rect 130 532 196 539
rect 327 582 414 649
rect 327 548 353 582
rect 387 548 414 582
rect 327 532 414 548
rect 647 560 751 572
rect 23 490 39 524
rect 73 498 89 524
rect 647 526 663 560
rect 697 526 751 560
rect 73 490 529 498
rect 23 464 529 490
rect 23 440 155 464
rect 23 406 39 440
rect 73 406 155 440
rect 23 390 155 406
rect 21 310 87 356
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 121 226 155 390
rect 37 192 155 226
rect 213 414 359 430
rect 213 380 236 414
rect 270 380 359 414
rect 213 364 359 380
rect 213 226 247 364
rect 281 310 359 326
rect 281 276 297 310
rect 331 276 359 310
rect 281 260 359 276
rect 395 320 461 430
rect 495 424 529 464
rect 647 492 751 526
rect 647 458 663 492
rect 697 458 751 492
rect 495 390 683 424
rect 395 286 411 320
rect 445 286 461 320
rect 395 270 461 286
rect 503 320 569 356
rect 503 286 519 320
rect 553 286 569 320
rect 503 270 569 286
rect 617 320 683 390
rect 617 286 633 320
rect 667 286 683 320
rect 617 270 683 286
rect 325 236 359 260
rect 717 236 751 458
rect 213 210 291 226
rect 213 192 241 210
rect 37 184 121 192
rect 37 150 53 184
rect 87 150 121 184
rect 225 176 241 192
rect 275 176 291 210
rect 325 210 751 236
rect 325 202 486 210
rect 37 108 121 150
rect 155 131 189 158
rect 155 17 189 97
rect 225 120 291 176
rect 470 176 486 202
rect 520 202 686 210
rect 520 176 536 202
rect 225 86 241 120
rect 275 86 291 120
rect 225 70 291 86
rect 325 147 427 156
rect 325 113 363 147
rect 397 113 427 147
rect 325 17 427 113
rect 470 140 536 176
rect 670 176 686 202
rect 720 176 751 210
rect 470 106 486 140
rect 520 106 536 140
rect 470 90 536 106
rect 570 146 636 168
rect 570 112 586 146
rect 620 112 636 146
rect 570 17 636 112
rect 670 140 751 176
rect 670 106 686 140
rect 720 106 751 140
rect 670 90 751 106
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or3b_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C_N
rlabel comment s 0 0 0 0 4 or3b_2
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 384 641 384 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 240 407 240 407 0 FreeSans 340 0 0 0 X
flabel locali s 336 407 336 407 0 FreeSans 340 0 0 0 X
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 A
flabel locali s 432 407 432 407 0 FreeSans 340 0 0 0 A
flabel locali s 528 333 528 333 0 FreeSans 340 0 0 0 B
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 C_N
rlabel comment s 0 0 0 0 4 or3b_2
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 384 641 384 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 240 407 240 407 0 FreeSans 340 0 0 0 X
flabel locali s 336 407 336 407 0 FreeSans 340 0 0 0 X
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 A
flabel locali s 432 407 432 407 0 FreeSans 340 0 0 0 A
flabel locali s 528 333 528 333 0 FreeSans 340 0 0 0 B
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 C_N
<< properties >>
string FIXED_BBOX 0 0 768 666
<< end >>
