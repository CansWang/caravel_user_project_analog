magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal1 >>
rect -195 -26 -186 26
rect -134 -26 -122 26
rect -70 -26 -58 26
rect -6 -26 6 26
rect 58 -26 70 26
rect 122 -26 134 26
rect 186 -26 195 26
<< via1 >>
rect -186 -26 -134 26
rect -122 -26 -70 26
rect -58 -26 -6 26
rect 6 -26 58 26
rect 70 -26 122 26
rect 134 -26 186 26
<< metal2 >>
rect -195 -26 -186 26
rect -134 -26 -122 26
rect -70 -26 -58 26
rect -6 -26 6 26
rect 58 -26 70 26
rect 122 -26 134 26
rect 186 -26 195 26
<< end >>
