magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< error_s >>
rect 542 31823 543 31868
rect 1790 31823 1791 31868
rect 3038 31823 3039 31868
rect 4958 31823 4959 31868
rect 6014 31823 6015 31868
rect 8126 31823 8127 31868
rect 9470 31823 9471 31868
rect 10334 31823 10335 31868
rect 12062 31823 12063 31868
rect 15902 31823 15903 31868
rect 17054 31823 17055 31868
rect 18494 31823 18495 31868
rect 19742 31823 19743 31868
rect 20990 31823 20991 31868
rect 22046 31823 22047 31868
rect 22910 31823 22911 31868
rect 24254 31823 24255 31868
rect 25502 31823 25503 31868
rect 26846 31823 26847 31868
rect 28094 31823 28095 31868
rect 29342 31823 29343 31868
rect 30686 31823 30687 31868
rect 1118 30747 1119 30792
rect 5630 30747 5631 30792
rect 7550 30747 7551 30792
rect 8798 30747 8799 30792
rect 10814 30747 10815 30792
rect 12062 30747 12063 30792
rect 13310 30747 13311 30792
rect 14558 30747 14559 30792
rect 15902 30747 15903 30792
rect 17150 30747 17151 30792
rect 18494 30747 18495 30792
rect 19550 30747 19551 30792
rect 20414 30747 20415 30792
rect 21662 30747 21663 30792
rect 22910 30747 22911 30792
rect 24254 30747 24255 30792
rect 25502 30747 25503 30792
rect 26846 30747 26847 30792
rect 28094 30747 28095 30792
rect 29342 30747 29343 30792
rect 30686 30747 30687 30792
rect 31550 30747 31551 30792
rect 542 30491 543 30536
rect 1790 30491 1791 30536
rect 6302 30491 6303 30536
rect 7070 30491 7071 30536
rect 8798 30491 8799 30536
rect 10814 30491 10815 30536
rect 12062 30491 12063 30536
rect 13310 30491 13311 30536
rect 14366 30491 14367 30536
rect 18494 30491 18495 30536
rect 19742 30491 19743 30536
rect 20990 30491 20991 30536
rect 22046 30491 22047 30536
rect 22910 30491 22911 30536
rect 24254 30491 24255 30536
rect 25502 30491 25503 30536
rect 26846 30491 26847 30536
rect 28094 30491 28095 30536
rect 29342 30491 29343 30536
rect 30686 30491 30687 30536
rect 1118 29415 1119 29460
rect 5630 29415 5631 29460
rect 6878 29415 6879 29460
rect 10814 29415 10815 29460
rect 15902 29415 15903 29460
rect 17150 29415 17151 29460
rect 18494 29415 18495 29460
rect 19550 29415 19551 29460
rect 20414 29415 20415 29460
rect 21662 29415 21663 29460
rect 22910 29415 22911 29460
rect 24254 29415 24255 29460
rect 25502 29415 25503 29460
rect 26846 29415 26847 29460
rect 28094 29415 28095 29460
rect 29342 29415 29343 29460
rect 30686 29415 30687 29460
rect 31550 29415 31551 29460
rect 542 29159 543 29204
rect 1790 29159 1791 29204
rect 3038 29159 3039 29204
rect 4382 29159 4383 29204
rect 5630 29159 5631 29204
rect 6878 29159 6879 29204
rect 9470 29159 9471 29204
rect 10814 29159 10815 29204
rect 13310 29159 13311 29204
rect 14654 29159 14655 29204
rect 15902 29159 15903 29204
rect 18494 29159 18495 29204
rect 19742 29159 19743 29204
rect 20990 29159 20991 29204
rect 22046 29159 22047 29204
rect 22910 29159 22911 29204
rect 24254 29159 24255 29204
rect 25502 29159 25503 29204
rect 26846 29159 26847 29204
rect 28094 29159 28095 29204
rect 29342 29159 29343 29204
rect 30686 29159 30687 29204
rect 1118 28083 1119 28128
rect 2462 28083 2463 28128
rect 3710 28083 3711 28128
rect 5534 28083 5535 28128
rect 6878 28083 6879 28128
rect 8222 28083 8223 28128
rect 9086 28083 9087 28128
rect 10814 28083 10815 28128
rect 11870 28083 11871 28128
rect 15902 28083 15903 28128
rect 17150 28083 17151 28128
rect 18494 28083 18495 28128
rect 19550 28083 19551 28128
rect 21662 28083 21663 28128
rect 22910 28083 22911 28128
rect 24254 28083 24255 28128
rect 28766 28083 28767 28128
rect 29534 28083 29535 28128
rect 30686 28083 30687 28128
rect 31550 28083 31551 28128
rect 542 27827 543 27872
rect 1790 27827 1791 27872
rect 3710 27827 3711 27872
rect 5630 27827 5631 27872
rect 10718 27827 10719 27872
rect 12062 27827 12063 27872
rect 13118 27827 13119 27872
rect 18494 27827 18495 27872
rect 19742 27827 19743 27872
rect 20990 27827 20991 27872
rect 22046 27827 22047 27872
rect 24254 27827 24255 27872
rect 27998 27827 27999 27872
rect 29342 27827 29343 27872
rect 30686 27827 30687 27872
rect 734 26751 735 26796
rect 8798 26751 8799 26796
rect 10814 26751 10815 26796
rect 12734 26751 12735 26796
rect 13982 26751 13983 26796
rect 15902 26751 15903 26796
rect 17150 26751 17151 26796
rect 18494 26751 18495 26796
rect 19550 26751 19551 26796
rect 21662 26751 21663 26796
rect 22910 26751 22911 26796
rect 24254 26751 24255 26796
rect 25502 26751 25503 26796
rect 26846 26751 26847 26796
rect 28094 26751 28095 26796
rect 29342 26751 29343 26796
rect 30686 26751 30687 26796
rect 31550 26751 31551 26796
rect 542 26495 543 26540
rect 1790 26495 1791 26540
rect 3038 26495 3039 26540
rect 4958 26495 4959 26540
rect 11390 26495 11391 26540
rect 12926 26495 12927 26540
rect 13982 26495 13983 26540
rect 15230 26495 15231 26540
rect 17054 26495 17055 26540
rect 20414 26495 20415 26540
rect 21662 26495 21663 26540
rect 25502 26495 25503 26540
rect 26846 26495 26847 26540
rect 30014 26495 30015 26540
rect 31262 26495 31263 26540
rect 4382 25419 4383 25464
rect 5630 25419 5631 25464
rect 15902 25419 15903 25464
rect 17150 25419 17151 25464
rect 19070 25419 19071 25464
rect 22334 25419 22335 25464
rect 23582 25419 23583 25464
rect 24542 25419 24543 25464
rect 28766 25419 28767 25464
rect 29534 25419 29535 25464
rect 30686 25419 30687 25464
rect 31550 25419 31551 25464
rect 542 25163 543 25208
rect 1790 25163 1791 25208
rect 3710 25163 3711 25208
rect 5534 25163 5535 25208
rect 6878 25163 6879 25208
rect 9470 25163 9471 25208
rect 11390 25163 11391 25208
rect 13310 25163 13311 25208
rect 15230 25163 15231 25208
rect 16094 25163 16095 25208
rect 18494 25163 18495 25208
rect 19358 25163 19359 25208
rect 22910 25163 22911 25208
rect 24254 25163 24255 25208
rect 25502 25163 25503 25208
rect 27038 25163 27039 25208
rect 28094 25163 28095 25208
rect 29342 25163 29343 25208
rect 31262 25163 31263 25208
rect 830 24087 831 24132
rect 2462 24087 2463 24132
rect 3710 24087 3711 24132
rect 6302 24087 6303 24132
rect 10814 24087 10815 24132
rect 12542 24087 12543 24132
rect 13790 24087 13791 24132
rect 16574 24087 16575 24132
rect 17822 24087 17823 24132
rect 19070 24087 19071 24132
rect 28094 24087 28095 24132
rect 29342 24087 29343 24132
rect 30686 24087 30687 24132
rect 31550 24087 31551 24132
rect 542 23831 543 23876
rect 1790 23831 1791 23876
rect 3710 23831 3711 23876
rect 4958 23831 4959 23876
rect 6206 23831 6207 23876
rect 8030 23831 8031 23876
rect 9374 23831 9375 23876
rect 10814 23831 10815 23876
rect 15902 23831 15903 23876
rect 18494 23831 18495 23876
rect 19742 23831 19743 23876
rect 20990 23831 20991 23876
rect 22046 23831 22047 23876
rect 22910 23831 22911 23876
rect 24254 23831 24255 23876
rect 25502 23831 25503 23876
rect 26846 23831 26847 23876
rect 28094 23831 28095 23876
rect 29342 23831 29343 23876
rect 31262 23831 31263 23876
rect 3806 22755 3807 22800
rect 6302 22755 6303 22800
rect 7550 22755 7551 22800
rect 8798 22755 8799 22800
rect 9566 22755 9567 22800
rect 10814 22755 10815 22800
rect 12062 22755 12063 22800
rect 13310 22755 13311 22800
rect 18398 22755 18399 22800
rect 20414 22755 20415 22800
rect 21662 22755 21663 22800
rect 23582 22755 23583 22800
rect 25502 22755 25503 22800
rect 26846 22755 26847 22800
rect 29342 22755 29343 22800
rect 30686 22755 30687 22800
rect 31550 22755 31551 22800
rect 542 22499 543 22544
rect 1790 22499 1791 22544
rect 4382 22499 4383 22544
rect 5150 22499 5151 22544
rect 6878 22499 6879 22544
rect 13310 22499 13311 22544
rect 14366 22499 14367 22544
rect 18494 22499 18495 22544
rect 24830 22499 24831 22544
rect 28094 22499 28095 22544
rect 30014 22499 30015 22544
rect 31262 22499 31263 22544
rect 3710 21423 3711 21468
rect 8798 21423 8799 21468
rect 9566 21423 9567 21468
rect 11102 21423 11103 21468
rect 12350 21423 12351 21468
rect 13598 21423 13599 21468
rect 15902 21423 15903 21468
rect 17630 21423 17631 21468
rect 22334 21423 22335 21468
rect 24254 21423 24255 21468
rect 28094 21423 28095 21468
rect 30686 21423 30687 21468
rect 31550 21423 31551 21468
rect 542 21167 543 21212
rect 1790 21167 1791 21212
rect 3710 21167 3711 21212
rect 4958 21167 4959 21212
rect 6206 21167 6207 21212
rect 11294 21167 11295 21212
rect 13982 21167 13983 21212
rect 15902 21167 15903 21212
rect 17054 21167 17055 21212
rect 20894 21167 20895 21212
rect 22046 21167 22047 21212
rect 25502 21167 25503 21212
rect 26846 21167 26847 21212
rect 29918 21167 29919 21212
rect 734 20091 735 20136
rect 2462 20091 2463 20136
rect 3614 20091 3615 20136
rect 10814 20091 10815 20136
rect 11870 20091 11871 20136
rect 15902 20091 15903 20136
rect 23582 20091 23583 20136
rect 24542 20091 24543 20136
rect 25502 20091 25503 20136
rect 26846 20091 26847 20136
rect 28094 20091 28095 20136
rect 29342 20091 29343 20136
rect 30686 20091 30687 20136
rect 31550 20091 31551 20136
rect 542 19835 543 19880
rect 1790 19835 1791 19880
rect 4958 19835 4959 19880
rect 6302 19835 6303 19880
rect 8222 19835 8223 19880
rect 13118 19835 13119 19880
rect 14270 19835 14271 19880
rect 18494 19835 18495 19880
rect 19742 19835 19743 19880
rect 20990 19835 20991 19880
rect 22046 19835 22047 19880
rect 22910 19835 22911 19880
rect 24350 19835 24351 19880
rect 28094 19835 28095 19880
rect 29342 19835 29343 19880
rect 3710 18759 3711 18804
rect 4574 18759 4575 18804
rect 5630 18759 5631 18804
rect 6878 18759 6879 18804
rect 8222 18759 8223 18804
rect 9470 18759 9471 18804
rect 10814 18759 10815 18804
rect 11582 18759 11583 18804
rect 13310 18759 13311 18804
rect 14558 18759 14559 18804
rect 15422 18759 15423 18804
rect 17150 18759 17151 18804
rect 22910 18759 22911 18804
rect 24254 18759 24255 18804
rect 30686 18759 30687 18804
rect 31550 18759 31551 18804
rect 542 18503 543 18548
rect 1790 18503 1791 18548
rect 3710 18503 3711 18548
rect 4958 18503 4959 18548
rect 6878 18503 6879 18548
rect 8606 18503 8607 18548
rect 10526 18503 10527 18548
rect 12062 18503 12063 18548
rect 13310 18503 13311 18548
rect 15230 18503 15231 18548
rect 16478 18503 16479 18548
rect 22910 18503 22911 18548
rect 24254 18503 24255 18548
rect 27998 18503 27999 18548
rect 29342 18503 29343 18548
rect 31262 18503 31263 18548
rect 5438 17427 5439 17472
rect 9470 17427 9471 17472
rect 11390 17427 11391 17472
rect 17438 17427 17439 17472
rect 21278 17427 21279 17472
rect 25406 17427 25407 17472
rect 26750 17427 26751 17472
rect 30686 17427 30687 17472
rect 31550 17427 31551 17472
rect 542 17171 543 17216
rect 1790 17171 1791 17216
rect 3902 17171 3903 17216
rect 4958 17171 4959 17216
rect 12062 17171 12063 17216
rect 20798 17171 20799 17216
rect 22046 17171 22047 17216
rect 30494 17171 30495 17216
rect 19550 16095 19551 16140
rect 20894 16095 20895 16140
rect 22334 16095 22335 16140
rect 24542 16095 24543 16140
rect 25502 16095 25503 16140
rect 27422 16095 27423 16140
rect 28766 16095 28767 16140
rect 29534 16095 29535 16140
rect 30686 16095 30687 16140
rect 31550 16095 31551 16140
rect 542 15839 543 15884
rect 1790 15839 1791 15884
rect 10814 15839 10815 15884
rect 12062 15839 12063 15884
rect 22910 15839 22911 15884
rect 24254 15839 24255 15884
rect 25502 15839 25503 15884
rect 26846 15839 26847 15884
rect 29342 15839 29343 15884
rect 31262 15839 31263 15884
rect 5630 14763 5631 14808
rect 6878 14763 6879 14808
rect 8222 14763 8223 14808
rect 9470 14763 9471 14808
rect 10814 14763 10815 14808
rect 12062 14763 12063 14808
rect 17150 14763 17151 14808
rect 18494 14763 18495 14808
rect 19550 14763 19551 14808
rect 20414 14763 20415 14808
rect 21662 14763 21663 14808
rect 28094 14763 28095 14808
rect 29342 14763 29343 14808
rect 30686 14763 30687 14808
rect 31550 14763 31551 14808
rect 542 14507 543 14552
rect 1790 14507 1791 14552
rect 3038 14507 3039 14552
rect 4382 14507 4383 14552
rect 10334 14507 10335 14552
rect 13886 14507 13887 14552
rect 15230 14507 15231 14552
rect 16574 14507 16575 14552
rect 20414 14507 20415 14552
rect 24254 14507 24255 14552
rect 25118 14507 25119 14552
rect 26846 14507 26847 14552
rect 30686 14507 30687 14552
rect 3902 13431 3903 13476
rect 12734 13431 12735 13476
rect 13982 13431 13983 13476
rect 15710 13431 15711 13476
rect 17150 13431 17151 13476
rect 18494 13431 18495 13476
rect 23582 13431 23583 13476
rect 26846 13431 26847 13476
rect 30686 13431 30687 13476
rect 31550 13431 31551 13476
rect 542 13175 543 13220
rect 1790 13175 1791 13220
rect 3038 13175 3039 13220
rect 14654 13175 14655 13220
rect 15902 13175 15903 13220
rect 17918 13175 17919 13220
rect 19646 13175 19647 13220
rect 25502 13175 25503 13220
rect 27038 13175 27039 13220
rect 30686 13175 30687 13220
rect 10622 12099 10623 12144
rect 13982 12099 13983 12144
rect 23582 12099 23583 12144
rect 26366 12099 26367 12144
rect 28094 12099 28095 12144
rect 30686 12099 30687 12144
rect 31550 12099 31551 12144
rect 1790 11843 1791 11888
rect 8222 11843 8223 11888
rect 9470 11843 9471 11888
rect 11390 11843 11391 11888
rect 12926 11843 12927 11888
rect 14462 11843 14463 11888
rect 18494 11843 18495 11888
rect 19742 11843 19743 11888
rect 22910 11843 22911 11888
rect 24254 11843 24255 11888
rect 25502 11843 25503 11888
rect 26846 11843 26847 11888
rect 28766 11843 28767 11888
rect 30014 11843 30015 11888
rect 31262 11843 31263 11888
rect 1790 10767 1791 10812
rect 2654 10767 2655 10812
rect 5630 10767 5631 10812
rect 6878 10767 6879 10812
rect 7646 10767 7647 10812
rect 10814 10767 10815 10812
rect 13694 10767 13695 10812
rect 16574 10767 16575 10812
rect 21662 10767 21663 10812
rect 22622 10767 22623 10812
rect 25502 10767 25503 10812
rect 26846 10767 26847 10812
rect 28094 10767 28095 10812
rect 29342 10767 29343 10812
rect 30686 10767 30687 10812
rect 31550 10767 31551 10812
rect 542 10511 543 10556
rect 3710 10511 3711 10556
rect 18398 10511 18399 10556
rect 19742 10511 19743 10556
rect 20990 10511 20991 10556
rect 22910 10511 22911 10556
rect 24830 10511 24831 10556
rect 26846 10511 26847 10556
rect 30686 10511 30687 10556
rect 926 9435 927 9480
rect 3326 9435 3327 9480
rect 4574 9435 4575 9480
rect 10814 9435 10815 9480
rect 12062 9435 12063 9480
rect 13982 9435 13983 9480
rect 15902 9435 15903 9480
rect 17150 9435 17151 9480
rect 18878 9435 18879 9480
rect 21374 9435 21375 9480
rect 22910 9435 22911 9480
rect 24254 9435 24255 9480
rect 28670 9435 28671 9480
rect 30686 9435 30687 9480
rect 31550 9435 31551 9480
rect 1502 9179 1503 9224
rect 5630 9179 5631 9224
rect 13310 9179 13311 9224
rect 15902 9179 15903 9224
rect 22910 9179 22911 9224
rect 24254 9179 24255 9224
rect 26174 9179 26175 9224
rect 28094 9179 28095 9224
rect 29342 9179 29343 9224
rect 30686 9179 30687 9224
rect 1022 8103 1023 8148
rect 5630 8103 5631 8148
rect 7262 8103 7263 8148
rect 9566 8103 9567 8148
rect 10814 8103 10815 8148
rect 12062 8103 12063 8148
rect 13982 8103 13983 8148
rect 15806 8103 15807 8148
rect 17150 8103 17151 8148
rect 18686 8103 18687 8148
rect 21374 8103 21375 8148
rect 22814 8103 22815 8148
rect 26846 8103 26847 8148
rect 27998 8103 27999 8148
rect 29342 8103 29343 8148
rect 30686 8103 30687 8148
rect 31550 8103 31551 8148
rect 542 7847 543 7892
rect 2078 7847 2079 7892
rect 3710 7847 3711 7892
rect 5630 7847 5631 7892
rect 6686 7847 6687 7892
rect 8222 7847 8223 7892
rect 9374 7847 9375 7892
rect 14654 7847 14655 7892
rect 17054 7847 17055 7892
rect 18494 7847 18495 7892
rect 19742 7847 19743 7892
rect 20990 7847 20991 7892
rect 22910 7847 22911 7892
rect 24254 7847 24255 7892
rect 25502 7847 25503 7892
rect 26846 7847 26847 7892
rect 28094 7847 28095 7892
rect 29342 7847 29343 7892
rect 30686 7847 30687 7892
rect 3038 6771 3039 6816
rect 4574 6771 4575 6816
rect 6782 6771 6783 6816
rect 13598 6771 13599 6816
rect 15710 6771 15711 6816
rect 16958 6771 16959 6816
rect 18302 6771 18303 6816
rect 20414 6771 20415 6816
rect 21662 6771 21663 6816
rect 22526 6771 22527 6816
rect 23774 6771 23775 6816
rect 28094 6771 28095 6816
rect 29342 6771 29343 6816
rect 30686 6771 30687 6816
rect 31550 6771 31551 6816
rect 542 6515 543 6560
rect 1790 6515 1791 6560
rect 3902 6515 3903 6560
rect 5438 6515 5439 6560
rect 13022 6515 13023 6560
rect 16574 6515 16575 6560
rect 21374 6515 21375 6560
rect 28094 6515 28095 6560
rect 29342 6515 29343 6560
rect 30686 6515 30687 6560
rect 11006 5439 11007 5484
rect 12542 5439 12543 5484
rect 15806 5439 15807 5484
rect 17150 5439 17151 5484
rect 25502 5439 25503 5484
rect 27422 5439 27423 5484
rect 28766 5439 28767 5484
rect 29534 5439 29535 5484
rect 30686 5439 30687 5484
rect 31550 5439 31551 5484
rect 542 5183 543 5228
rect 1790 5183 1791 5228
rect 6494 5183 6495 5228
rect 9182 5183 9183 5228
rect 10430 5183 10431 5228
rect 14654 5183 14655 5228
rect 18494 5183 18495 5228
rect 20414 5183 20415 5228
rect 22046 5183 22047 5228
rect 25502 5183 25503 5228
rect 26846 5183 26847 5228
rect 30686 5183 30687 5228
rect 4382 4107 4383 4152
rect 5630 4107 5631 4152
rect 6878 4107 6879 4152
rect 8222 4107 8223 4152
rect 12734 4107 12735 4152
rect 13886 4107 13887 4152
rect 16190 4107 16191 4152
rect 17342 4107 17343 4152
rect 18590 4107 18591 4152
rect 22910 4107 22911 4152
rect 23774 4107 23775 4152
rect 25502 4107 25503 4152
rect 27806 4107 27807 4152
rect 29342 4107 29343 4152
rect 30686 4107 30687 4152
rect 31550 4107 31551 4152
rect 542 3851 543 3896
rect 1790 3851 1791 3896
rect 3710 3851 3711 3896
rect 5342 3851 5343 3896
rect 6878 3851 6879 3896
rect 10142 3851 10143 3896
rect 11390 3851 11391 3896
rect 13310 3851 13311 3896
rect 14270 3851 14271 3896
rect 19070 3851 19071 3896
rect 23582 3851 23583 3896
rect 24830 3851 24831 3896
rect 26846 3851 26847 3896
rect 28094 3851 28095 3896
rect 29342 3851 29343 3896
rect 30686 3851 30687 3896
rect 1118 2775 1119 2820
rect 2462 2775 2463 2820
rect 3710 2775 3711 2820
rect 6110 2775 6111 2820
rect 7550 2775 7551 2820
rect 8510 2775 8511 2820
rect 9566 2775 9567 2820
rect 12062 2775 12063 2820
rect 13982 2775 13983 2820
rect 15902 2775 15903 2820
rect 17342 2775 17343 2820
rect 20414 2775 20415 2820
rect 22334 2775 22335 2820
rect 23582 2775 23583 2820
rect 25502 2775 25503 2820
rect 26846 2775 26847 2820
rect 30686 2775 30687 2820
rect 31550 2775 31551 2820
rect 542 2519 543 2564
rect 1790 2519 1791 2564
rect 3998 2519 3999 2564
rect 6878 2519 6879 2564
rect 7934 2519 7935 2564
rect 9470 2519 9471 2564
rect 11390 2519 11391 2564
rect 18494 2519 18495 2564
rect 19550 2519 19551 2564
rect 22910 2519 22911 2564
rect 24254 2519 24255 2564
rect 28094 2519 28095 2564
rect 29342 2519 29343 2564
rect 30686 2519 30687 2564
rect 1118 1443 1119 1488
rect 2270 1443 2271 1488
rect 4382 1443 4383 1488
rect 9566 1443 9567 1488
rect 13310 1443 13311 1488
rect 15902 1443 15903 1488
rect 17150 1443 17151 1488
rect 18494 1443 18495 1488
rect 19550 1443 19551 1488
rect 20414 1443 20415 1488
rect 21662 1443 21663 1488
rect 22910 1443 22911 1488
rect 25502 1443 25503 1488
rect 26846 1443 26847 1488
rect 28094 1443 28095 1488
rect 29342 1443 29343 1488
rect 30686 1443 30687 1488
rect 31550 1443 31551 1488
rect 542 1187 543 1232
rect 1790 1187 1791 1232
rect 5630 1187 5631 1232
rect 6878 1187 6879 1232
rect 8222 1187 8223 1232
rect 9470 1187 9471 1232
rect 10814 1187 10815 1232
rect 12062 1187 12063 1232
rect 13982 1187 13983 1232
rect 15230 1187 15231 1232
rect 16574 1187 16575 1232
rect 19070 1187 19071 1232
rect 20414 1187 20415 1232
rect 21662 1187 21663 1232
rect 22910 1187 22911 1232
rect 24254 1187 24255 1232
rect 25502 1187 25503 1232
rect 26846 1187 26847 1232
rect 28094 1187 28095 1232
rect 29342 1187 29343 1232
rect 30686 1187 30687 1232
rect 1118 111 1119 156
rect 2078 111 2079 156
rect 3038 111 3039 156
rect 4382 111 4383 156
rect 5630 111 5631 156
rect 6878 111 6879 156
rect 8222 111 8223 156
rect 9470 111 9471 156
rect 10814 111 10815 156
rect 12062 111 12063 156
rect 13310 111 13311 156
rect 14558 111 14559 156
rect 15902 111 15903 156
rect 17054 111 17055 156
rect 18494 111 18495 156
rect 19550 111 19551 156
rect 20414 111 20415 156
rect 21662 111 21663 156
rect 22910 111 22911 156
rect 24254 111 24255 156
rect 25502 111 25503 156
rect 26846 111 26847 156
rect 28094 111 28095 156
rect 29342 111 29343 156
rect 30686 111 30687 156
<< locali >>
rect 6367 31618 6480 31652
rect 6672 31618 6785 31652
rect 10687 31618 10800 31652
rect 11184 31618 11297 31652
rect 6367 31544 6401 31618
rect 6751 31396 6785 31618
rect 11263 31470 11297 31618
rect 8095 30360 8208 30394
rect 8095 30064 8129 30360
rect 16255 29546 16368 29580
rect 16255 29398 16289 29546
rect 16735 28988 16769 29136
rect 12031 28880 12065 28971
rect 12144 28954 12257 28988
rect 12223 28732 12257 28954
rect 16351 28954 16464 28988
rect 16656 28954 16769 28988
rect 16351 28732 16385 28954
rect 4752 28288 4865 28322
rect 4255 28214 4368 28248
rect 4831 28066 4865 28288
rect 6559 27730 6593 27878
rect 2815 27696 2928 27730
rect 3120 27696 3233 27730
rect 2815 27400 2849 27696
rect 3199 27400 3233 27696
rect 6175 27696 6288 27730
rect 6480 27696 6593 27730
rect 11071 27730 11105 27878
rect 11071 27696 11184 27730
rect 11376 27696 11489 27730
rect 4351 27582 4385 27639
rect 4848 27622 4961 27656
rect 4159 27548 4385 27582
rect 4159 27474 4193 27548
rect 4927 27400 4961 27622
rect 6175 27548 6209 27696
rect 11455 27400 11489 27696
rect 13471 27656 13505 27878
rect 23664 27696 23777 27730
rect 13471 27622 13584 27656
rect 13663 27400 13697 27639
rect 23743 27400 23777 27696
rect 1567 26973 1601 27212
rect 1680 26956 1793 26990
rect 1759 26734 1793 26956
rect 9631 26916 9665 27212
rect 9552 26882 9665 26916
rect 18559 26398 18593 26472
rect 18559 26364 18768 26398
rect 3967 26290 4080 26324
rect 5695 26290 5808 26324
rect 3967 26068 4001 26290
rect 5695 26068 5729 26290
rect 16159 26068 16193 26307
rect 6751 25658 6785 25880
rect 6672 25624 6785 25658
rect 7807 25584 7841 25880
rect 9631 25658 9665 25880
rect 9552 25624 9665 25658
rect 12223 25658 12257 25732
rect 12223 25624 12336 25658
rect 16639 25584 16673 25732
rect 7807 25550 8016 25584
rect 8304 25550 8417 25584
rect 8383 25402 8417 25550
rect 10879 25550 11184 25584
rect 16255 25550 16368 25584
rect 16560 25550 16673 25584
rect 10879 25476 10913 25550
rect 16255 25402 16289 25550
rect 4063 24992 4097 25214
rect 14047 25032 14160 25066
rect 26047 25032 26160 25066
rect 4063 24958 4176 24992
rect 10896 24958 11009 24992
rect 10975 24884 11009 24958
rect 11839 24884 12048 24918
rect 11839 24736 11873 24884
rect 14047 24736 14081 25032
rect 26047 24736 26081 25032
rect 11551 24252 11585 24548
rect 14527 24326 14561 24474
rect 14448 24292 14561 24326
rect 1584 24218 1697 24252
rect 11551 24218 11664 24252
rect 11856 24218 11969 24252
rect 1663 24070 1697 24218
rect 11935 24070 11969 24218
rect 2815 23660 2849 23882
rect 7248 23700 7361 23734
rect 2815 23626 2928 23660
rect 7327 23404 7361 23700
rect 9727 23660 9761 23882
rect 8383 23586 8417 23660
rect 9727 23626 9840 23660
rect 8383 23552 8496 23586
rect 9919 23404 9953 23643
rect 11359 23552 11393 23643
rect 4560 23182 4673 23216
rect 13663 22994 13697 23216
rect 4639 22920 4673 22994
rect 4159 22886 4272 22920
rect 4560 22886 4673 22920
rect 13663 22960 13776 22994
rect 27871 22960 27984 22994
rect 4159 22812 4193 22886
rect 13663 22738 13697 22960
rect 25855 22886 25968 22920
rect 25855 22738 25889 22886
rect 27871 22812 27905 22960
rect 3007 22328 3041 22550
rect 6271 22402 6305 22550
rect 6192 22368 6305 22402
rect 8863 22368 9072 22402
rect 23376 22368 23760 22402
rect 3007 22294 3120 22328
rect 3199 22072 3233 22311
rect 8016 22294 8225 22328
rect 8191 22220 8225 22294
rect 25584 22220 25793 22254
rect 5791 21662 5825 21736
rect 5712 21628 5825 21662
rect 7903 21662 7937 21884
rect 7903 21628 8016 21662
rect 14335 21588 14369 21884
rect 16447 21662 16481 21810
rect 16447 21628 16560 21662
rect 16639 21645 16673 21884
rect 19920 21628 20112 21662
rect 13951 21554 14064 21588
rect 14256 21554 14369 21588
rect 18751 21554 18864 21588
rect 13951 21406 13985 21554
rect 18751 21480 18785 21554
rect 28543 21440 28577 21810
rect 28543 21406 28656 21440
rect 5407 21070 5441 21218
rect 11647 21070 11681 21218
rect 4063 21036 4176 21070
rect 5407 21036 5520 21070
rect 8592 21036 9456 21070
rect 11647 21036 11760 21070
rect 5407 20740 5441 21036
rect 6559 20962 6672 20996
rect 6559 20740 6593 20962
rect 7135 20888 7169 20979
rect 9055 20740 9089 21036
rect 10303 20962 10416 20996
rect 30271 20962 30384 20996
rect 10303 20740 10337 20962
rect 30271 20740 30305 20962
rect 1567 20313 1601 20552
rect 4560 20296 4673 20330
rect 5503 20256 5537 20330
rect 3967 20222 4080 20256
rect 5503 20222 5712 20256
rect 3967 20148 4001 20222
rect 6751 19704 6864 19738
rect 4464 19630 4577 19664
rect 4543 19556 4577 19630
rect 6751 19556 6785 19704
rect 9264 19630 9377 19664
rect 13471 19630 13584 19664
rect 13776 19630 13889 19664
rect 13471 19408 13505 19630
rect 13855 19482 13889 19630
rect 15967 18981 16001 19072
rect 17503 18890 17616 18924
rect 17503 18742 17537 18890
rect 3295 18332 3329 18554
rect 10879 18372 10992 18406
rect 3216 18298 3329 18332
rect 5695 18224 5729 18315
rect 6192 18298 6305 18332
rect 6271 18150 6305 18298
rect 10879 18224 10913 18372
rect 17023 18076 17057 18315
rect 7248 17854 7361 17888
rect 16447 17706 16752 17740
rect 6096 17632 6497 17666
rect 6463 17592 6497 17632
rect 7999 17592 8033 17649
rect 6463 17558 6864 17592
rect 7903 17558 8033 17592
rect 12703 17632 12816 17666
rect 13200 17632 13313 17666
rect 6655 17484 6689 17558
rect 7903 17410 7937 17558
rect 12703 17484 12737 17632
rect 16447 17592 16481 17706
rect 15792 17558 16481 17592
rect 16639 17558 16673 17706
rect 19807 17666 19841 17814
rect 18271 17632 18672 17666
rect 19728 17632 19841 17666
rect 18271 17592 18305 17632
rect 18096 17558 18305 17592
rect 25759 17558 25872 17592
rect 18175 17410 18209 17558
rect 25759 17410 25793 17558
rect 3007 17074 3041 17148
rect 3007 17040 3120 17074
rect 3408 17040 3521 17074
rect 5311 17000 5345 17148
rect 8863 17000 8897 17148
rect 9247 17000 9281 17222
rect 10687 17000 10721 17222
rect 11647 17074 11681 17222
rect 11568 17040 11681 17074
rect 5311 16966 5424 17000
rect 8479 16818 8513 16983
rect 8863 16966 8976 17000
rect 9168 16966 9281 17000
rect 9840 16966 9953 17000
rect 10608 16966 10721 17000
rect 28639 16966 28752 17000
rect 9919 16744 9953 16966
rect 28639 16892 28673 16966
rect 9055 16260 9089 16556
rect 14047 16300 14160 16334
rect 14239 16317 14273 16408
rect 23359 16334 23393 16408
rect 25855 16334 25889 16556
rect 18768 16300 18881 16334
rect 23359 16300 23472 16334
rect 25855 16300 25968 16334
rect 8287 16226 8400 16260
rect 8592 16226 9264 16260
rect 8287 16152 8321 16226
rect 13567 16186 13601 16260
rect 13488 16152 13601 16186
rect 14047 16152 14081 16300
rect 18847 16078 18881 16300
rect 18480 15708 18593 15742
rect 18559 15412 18593 15708
rect 4063 14928 4097 15002
rect 4063 14894 4176 14928
rect 5983 14336 6017 14484
rect 7135 14410 7169 14558
rect 9535 14410 9569 14558
rect 7135 14376 7248 14410
rect 8575 14336 8609 14410
rect 9535 14376 9648 14410
rect 5983 14302 6096 14336
rect 8575 14302 8688 14336
rect 11551 14302 11664 14336
rect 11551 14080 11585 14302
rect 11743 14228 11777 14319
rect 14719 14080 14753 14319
rect 18096 14302 18209 14336
rect 26064 14302 26177 14336
rect 18175 14154 18209 14302
rect 26143 14080 26177 14302
rect 9840 13636 10224 13670
rect 11359 13596 11393 13892
rect 4752 13562 4865 13596
rect 11280 13562 11393 13596
rect 17791 13596 17825 13892
rect 21535 13670 21569 13818
rect 23167 13670 23201 13892
rect 21456 13636 21569 13670
rect 23088 13636 23201 13670
rect 24223 13596 24257 13744
rect 17791 13562 17904 13596
rect 19440 13562 19553 13596
rect 24223 13562 24336 13596
rect 19519 13414 19553 13562
rect 13855 13004 13889 13226
rect 15391 13078 15425 13226
rect 16831 13078 16865 13226
rect 15007 13044 15120 13078
rect 15312 13044 15425 13078
rect 16752 13044 16865 13078
rect 3696 12970 3792 13004
rect 5232 12970 5328 13004
rect 13855 12970 13968 13004
rect 14160 12970 14273 13004
rect 14239 12822 14273 12970
rect 15007 12896 15041 13044
rect 4464 12304 4577 12338
rect 4543 12230 4577 12304
rect 11359 12264 11393 12486
rect 14335 12338 14369 12560
rect 17023 12338 17057 12486
rect 14335 12304 14448 12338
rect 14640 12304 14753 12338
rect 16944 12304 17057 12338
rect 17503 12338 17537 12560
rect 17503 12304 17616 12338
rect 20767 12321 20801 12412
rect 11280 12230 11393 12264
rect 14719 12082 14753 12304
rect 23935 12264 23969 12412
rect 27216 12304 27329 12338
rect 29215 12321 29249 12412
rect 29328 12304 29441 12338
rect 23935 12230 24048 12264
rect 27295 12156 27329 12304
rect 29407 12156 29441 12304
rect 27871 11746 27905 11894
rect 8671 11712 8784 11746
rect 27871 11712 27984 11746
rect 8671 11564 8705 11712
rect 13471 11564 13505 11655
rect 20688 11638 20801 11672
rect 20767 11416 20801 11638
rect 4831 11006 4865 11228
rect 991 10972 1104 11006
rect 1296 10972 1409 11006
rect 4752 10972 4865 11006
rect 7999 11006 8033 11228
rect 8863 11006 8897 11228
rect 14047 11006 14081 11228
rect 18655 11006 18689 11228
rect 7999 10972 8112 11006
rect 8304 10972 9456 11006
rect 9840 10972 9953 11006
rect 14047 10972 14160 11006
rect 991 10750 1025 10972
rect 1375 10750 1409 10972
rect 9919 10750 9953 10972
rect 15679 10932 15713 11006
rect 18480 10972 18689 11006
rect 20287 10932 20321 11228
rect 24607 11006 24641 11228
rect 23472 10972 23585 11006
rect 24528 10972 24641 11006
rect 12703 10898 12912 10932
rect 13200 10898 13313 10932
rect 15679 10898 15792 10932
rect 19135 10898 19248 10932
rect 19536 10898 19649 10932
rect 20287 10898 20400 10932
rect 12703 10750 12737 10898
rect 19615 10750 19649 10898
rect 23551 10750 23585 10972
rect 26352 10898 26465 10932
rect 26431 10750 26465 10898
rect 13279 10414 13313 10562
rect 13200 10380 13313 10414
rect 21631 10414 21665 10488
rect 21631 10380 21744 10414
rect 25855 10340 25889 10562
rect 26239 10340 26273 10488
rect 11952 10306 12065 10340
rect 15984 10306 16368 10340
rect 22032 10306 22145 10340
rect 12031 10232 12065 10306
rect 22111 10232 22145 10306
rect 23551 10306 23664 10340
rect 25855 10306 25968 10340
rect 26160 10306 26273 10340
rect 10320 10084 10433 10118
rect 23551 10084 23585 10306
rect 1584 9640 1697 9674
rect 2335 9640 2448 9674
rect 1663 9418 1697 9640
rect 12511 9600 12545 9896
rect 17983 9640 18096 9674
rect 12511 9566 12624 9600
rect 17983 9418 18017 9640
rect 20863 9600 20897 9896
rect 21727 9674 21761 9748
rect 21727 9640 21840 9674
rect 20191 9566 20304 9600
rect 20784 9566 20897 9600
rect 23455 9600 23489 9896
rect 23455 9566 23568 9600
rect 20191 9418 20225 9566
rect 3967 8752 4001 9156
rect 5215 9008 5249 9156
rect 13855 9082 13889 9230
rect 13855 9048 14064 9082
rect 14352 9048 14945 9082
rect 19440 9048 19553 9082
rect 5136 8974 5249 9008
rect 13951 8752 13985 9048
rect 14911 9008 14945 9048
rect 14911 8974 15312 9008
rect 16351 8974 16560 9008
rect 16351 8826 16385 8974
rect 19519 8752 19553 9048
rect 21055 9008 21089 9230
rect 20784 8974 21089 9008
rect 24799 9008 24833 9230
rect 26928 9048 27041 9082
rect 24799 8974 24912 9008
rect 24991 8752 25025 8991
rect 27007 8752 27041 9048
rect 12799 8530 12912 8564
rect 1759 8268 1793 8416
rect 13087 8399 13121 8490
rect 1680 8234 1793 8268
rect 18192 8234 18305 8268
rect 20095 8120 20129 8490
rect 21727 8268 21761 8564
rect 24223 8268 24257 8490
rect 24607 8268 24641 8564
rect 25759 8325 25793 8564
rect 25951 8342 25985 8416
rect 25872 8308 25985 8342
rect 28351 8342 28385 8416
rect 28351 8308 28464 8342
rect 21727 8234 21840 8268
rect 22128 8234 22241 8268
rect 24223 8234 24336 8268
rect 24528 8234 24641 8268
rect 21727 8160 21761 8234
rect 20095 8086 20208 8120
rect 22207 8086 22241 8234
rect 1663 7750 1697 7898
rect 1584 7716 1697 7750
rect 10128 7716 10800 7750
rect 12048 7716 12161 7750
rect 10399 7420 10433 7716
rect 12127 7420 12161 7716
rect 15679 7676 15713 7898
rect 15487 7568 15521 7659
rect 15600 7642 15713 7676
rect 2431 6936 2465 7084
rect 5520 6976 5633 7010
rect 7440 6976 7553 7010
rect 2352 6902 2465 6936
rect 5599 6754 5633 6976
rect 7519 6754 7553 6976
rect 8479 6936 8513 7158
rect 14431 7010 14465 7232
rect 14352 6976 14465 7010
rect 17311 6936 17345 7010
rect 24127 6976 24240 7010
rect 8400 6902 8513 6936
rect 10704 6902 11088 6936
rect 17311 6902 17424 6936
rect 24127 6754 24161 6976
rect 3007 6344 3041 6566
rect 4255 6344 4289 6566
rect 13375 6418 13409 6566
rect 13375 6384 13488 6418
rect 23647 6344 23681 6418
rect 3007 6310 3120 6344
rect 4255 6310 4368 6344
rect 23568 6310 23681 6344
rect 25279 6344 25313 6418
rect 25279 6310 25392 6344
rect 25776 6310 26736 6344
rect 13200 5644 13313 5678
rect 14256 5644 15137 5678
rect 16639 5661 16673 5900
rect 11952 5570 12065 5604
rect 12031 5496 12065 5570
rect 13279 5496 13313 5644
rect 15103 5604 15137 5644
rect 15103 5570 15216 5604
rect 15103 5422 15137 5570
rect 10783 5086 10817 5160
rect 8287 5052 8400 5086
rect 9535 5052 9648 5086
rect 9840 5052 9953 5086
rect 10783 5052 10896 5086
rect 23184 5052 23681 5086
rect 7327 4904 7361 4995
rect 7440 4978 7649 5012
rect 7615 4830 7649 4978
rect 8287 4756 8321 5052
rect 9535 4904 9569 5052
rect 9919 4830 9953 5052
rect 23647 5012 23681 5052
rect 24223 5012 24257 5234
rect 20863 4938 20897 4995
rect 23647 4978 24336 5012
rect 20767 4904 20897 4938
rect 20767 4756 20801 4904
rect 1584 4312 1793 4346
rect 13183 4272 13217 4494
rect 26527 4272 26561 4420
rect 28639 4329 28673 4420
rect 912 4238 1025 4272
rect 13183 4238 13296 4272
rect 14239 4238 14352 4272
rect 20784 4238 20897 4272
rect 26448 4238 26561 4272
rect 14239 4090 14273 4238
rect 20863 4090 20897 4238
rect 4447 3720 4560 3754
rect 4447 3498 4481 3720
rect 18559 3680 18593 3902
rect 18480 3646 18593 3680
rect 22879 3680 22913 3828
rect 26143 3680 26177 3828
rect 22879 3646 22992 3680
rect 26064 3646 26177 3680
rect 5311 2940 5345 3162
rect 13087 2997 13121 3236
rect 22687 2940 22721 3162
rect 23167 2940 23201 3236
rect 24607 3014 24641 3236
rect 24528 2980 24641 3014
rect 5311 2906 5424 2940
rect 10687 2906 10800 2940
rect 22687 2906 22800 2940
rect 23088 2906 23201 2940
rect 10687 2758 10721 2906
rect 5599 2348 5633 2496
rect 5520 2314 5633 2348
rect 10495 2348 10529 2422
rect 10879 2348 10913 2570
rect 8767 2240 8801 2331
rect 10495 2314 10608 2348
rect 10800 2314 10913 2348
rect 14239 1648 14352 1682
rect 14431 1665 14465 1756
rect 14239 1426 14273 1648
rect 20767 1608 20801 1830
rect 23935 1665 23969 1756
rect 20767 1574 20880 1608
rect 13471 1090 13505 1238
rect 13392 1056 13505 1090
rect 17887 1056 18000 1090
rect 3600 982 3713 1016
rect 17887 834 17921 1056
<< metal1 >>
rect 0 32585 32064 32683
rect 34 32361 24734 32389
rect 24706 32287 24734 32361
rect 0 31919 32064 32017
rect 10690 31769 12638 31797
rect 10690 31649 10718 31769
rect 12610 31695 12638 31769
rect 2050 31621 4190 31649
rect 8578 31621 8702 31649
rect 8770 31621 10718 31649
rect 12322 31621 13022 31649
rect 4258 31547 6590 31575
rect 11458 31547 12158 31575
rect 11458 31501 11486 31547
rect 11266 31473 11486 31501
rect 12130 31501 12158 31547
rect 12130 31473 12734 31501
rect 12706 31464 12734 31473
rect 14626 31473 14846 31501
rect 14626 31464 14654 31473
rect 12706 31436 14654 31464
rect 6274 31399 6590 31427
rect 6681 31399 6768 31427
rect 8290 31399 8702 31427
rect 0 31253 32064 31351
rect 1977 31177 2064 31205
rect 30082 31177 30302 31205
rect 2530 31140 4190 31168
rect 2530 31131 2558 31140
rect 34 31103 254 31131
rect 226 31057 254 31103
rect 2338 31103 2558 31131
rect 4162 31131 4190 31140
rect 4162 31103 6974 31131
rect 226 31029 1886 31057
rect 1858 30983 1886 31029
rect 2338 30983 2366 31103
rect 6946 31057 6974 31103
rect 8194 31103 9758 31131
rect 8194 31057 8222 31103
rect 6946 31029 8222 31057
rect 9730 31057 9758 31103
rect 21634 31103 21854 31131
rect 21634 31057 21662 31103
rect 9730 31029 21662 31057
rect 21826 31029 21854 31103
rect 30274 31057 30302 31177
rect 31810 31177 32030 31205
rect 31810 31057 31838 31177
rect 30274 31029 31838 31057
rect 1858 30955 2366 30983
rect 3298 30955 3902 30983
rect 6562 30955 6686 30983
rect 8674 30955 9470 30983
rect 4258 30881 5918 30909
rect 6274 30881 6494 30909
rect 6681 30881 6768 30909
rect 8386 30881 9278 30909
rect 9465 30881 9552 30909
rect 5890 30835 5918 30881
rect 5890 30807 6590 30835
rect 7618 30807 8222 30835
rect 7618 30761 7646 30807
rect 8194 30798 8222 30807
rect 8194 30770 9182 30798
rect 7426 30733 7646 30761
rect 9154 30761 9182 30770
rect 9154 30733 9374 30761
rect 0 30587 32064 30685
rect 8674 30511 8894 30539
rect 8866 30465 8894 30511
rect 9346 30511 9566 30539
rect 9346 30465 9374 30511
rect 6754 30437 6974 30465
rect 6946 30391 6974 30437
rect 8002 30437 8222 30465
rect 8866 30437 9374 30465
rect 8002 30391 8030 30437
rect 6946 30363 8030 30391
rect 8290 30363 8414 30391
rect 13858 30363 15326 30391
rect 3225 30289 3312 30317
rect 9657 30289 9744 30317
rect 13858 30243 13886 30363
rect 2050 30215 2942 30243
rect 13474 30215 13886 30243
rect 15298 30243 15326 30363
rect 16953 30289 17040 30317
rect 17122 30289 17438 30317
rect 15298 30215 15696 30243
rect 14146 30141 15038 30169
rect 14146 30095 14174 30141
rect 4738 30067 5150 30095
rect 8098 30067 8510 30095
rect 13954 30067 14174 30095
rect 15010 30095 15038 30141
rect 15010 30067 15230 30095
rect 0 29921 32064 30019
rect 1954 29845 2078 29873
rect 9538 29845 9758 29873
rect 16642 29845 17150 29873
rect 2914 29808 5342 29836
rect 2914 29799 2942 29808
rect 2722 29771 2942 29799
rect 5314 29799 5342 29808
rect 12034 29808 13982 29836
rect 12034 29799 12062 29808
rect 5314 29771 5534 29799
rect 5698 29771 6302 29799
rect 11842 29771 12062 29799
rect 13954 29799 13982 29808
rect 13954 29771 14174 29799
rect 5698 29725 5726 29771
rect 3106 29697 3216 29725
rect 4834 29697 5726 29725
rect 6274 29725 6302 29771
rect 6274 29697 7166 29725
rect 7330 29697 7454 29725
rect 9072 29697 12144 29725
rect 4834 29651 4862 29697
rect 7138 29651 7166 29697
rect 2073 29623 2160 29651
rect 2722 29623 3614 29651
rect 3586 29614 3614 29623
rect 4354 29623 4862 29651
rect 4930 29623 5150 29651
rect 4354 29614 4382 29623
rect 3586 29586 4382 29614
rect 5122 29614 5150 29623
rect 5794 29623 6014 29651
rect 7138 29623 7742 29651
rect 12249 29623 12542 29651
rect 5794 29614 5822 29623
rect 5122 29586 5822 29614
rect 226 29549 1694 29577
rect 1881 29549 1968 29577
rect 2242 29549 3326 29577
rect 7522 29549 7550 29623
rect 12514 29614 12542 29623
rect 13762 29623 14558 29651
rect 16377 29623 16464 29651
rect 30946 29623 31934 29651
rect 13762 29614 13790 29623
rect 12514 29586 13790 29614
rect 11865 29549 11952 29577
rect 14722 29549 16190 29577
rect 16569 29549 16656 29577
rect 16834 29549 22142 29577
rect 226 29503 254 29549
rect 34 29475 254 29503
rect 1666 29503 1694 29549
rect 14722 29503 14750 29549
rect 1666 29475 1886 29503
rect 1858 29466 1886 29475
rect 3394 29475 14750 29503
rect 16162 29503 16190 29549
rect 16834 29503 16862 29549
rect 16162 29475 16862 29503
rect 22114 29503 22142 29549
rect 22114 29475 22334 29503
rect 3394 29466 3422 29475
rect 1858 29438 3422 29466
rect 16185 29401 16272 29429
rect 0 29255 32064 29353
rect 11650 29179 11966 29207
rect 14050 29105 16766 29133
rect 11458 29031 13982 29059
rect 6754 28957 8222 28985
rect 8290 28957 8414 28985
rect 8496 28957 8583 28985
rect 9826 28957 11870 28985
rect 13858 28957 13886 29031
rect 14146 28957 16190 28985
rect 14146 28911 14174 28957
rect 11961 28883 14174 28911
rect 16162 28911 16190 28957
rect 16162 28883 16670 28911
rect 14146 28772 16094 28800
rect 14146 28763 14174 28772
rect 7906 28735 8030 28763
rect 11842 28735 12254 28763
rect 13954 28735 14174 28763
rect 16066 28763 16094 28772
rect 16066 28735 16382 28763
rect 0 28589 32064 28687
rect 5913 28513 6000 28541
rect 13186 28476 14942 28504
rect 13186 28467 13214 28476
rect 130 28439 350 28467
rect 322 28393 350 28439
rect 1954 28439 4478 28467
rect 1954 28393 1982 28439
rect 322 28365 1982 28393
rect 4450 28393 4478 28439
rect 5314 28439 6878 28467
rect 5314 28393 5342 28439
rect 6850 28393 6878 28439
rect 9250 28439 10046 28467
rect 9250 28393 9278 28439
rect 4450 28365 5342 28393
rect 5506 28365 6494 28393
rect 6850 28365 9278 28393
rect 10018 28393 10046 28439
rect 12994 28439 13214 28467
rect 14914 28467 14942 28476
rect 14914 28439 15134 28467
rect 12994 28393 13022 28439
rect 10018 28365 13022 28393
rect 15106 28393 15134 28439
rect 18466 28439 21086 28467
rect 18466 28393 18494 28439
rect 15106 28365 18494 28393
rect 21058 28393 21086 28439
rect 23842 28439 24062 28467
rect 23842 28393 23870 28439
rect 21058 28365 23870 28393
rect 28066 28365 28478 28393
rect 2146 28291 3230 28319
rect 3312 28291 3399 28319
rect 6105 28291 6192 28319
rect 3202 28245 3230 28291
rect 6370 28245 6398 28319
rect 6466 28291 6494 28365
rect 9442 28291 9566 28319
rect 9730 28291 9854 28319
rect 14457 28291 14544 28319
rect 20674 28291 20894 28319
rect 25474 28291 26270 28319
rect 26242 28282 26270 28291
rect 27490 28291 27710 28319
rect 27490 28282 27518 28291
rect 26242 28254 27518 28282
rect 3202 28217 4286 28245
rect 6370 28217 6686 28245
rect 14050 28217 14942 28245
rect 18658 28217 20606 28245
rect 2338 28143 3038 28171
rect 2338 28097 2366 28143
rect 2146 28069 2366 28097
rect 3010 28097 3038 28143
rect 25954 28143 27518 28171
rect 25954 28097 25982 28143
rect 3010 28069 3230 28097
rect 4738 28069 4862 28097
rect 9250 28069 9662 28097
rect 12537 28069 12624 28097
rect 21058 28069 21182 28097
rect 25762 28069 25982 28097
rect 27490 28097 27518 28143
rect 27490 28069 27710 28097
rect 0 27923 32064 28021
rect 6178 27847 6302 27875
rect 6562 27847 6686 27875
rect 8674 27847 8894 27875
rect 8866 27838 8894 27847
rect 9730 27847 9950 27875
rect 11074 27847 11294 27875
rect 9730 27838 9758 27847
rect 8866 27810 9758 27838
rect 11266 27838 11294 27847
rect 11842 27847 12062 27875
rect 12610 27847 12830 27875
rect 11842 27838 11870 27847
rect 11266 27810 11870 27838
rect 12802 27801 12830 27847
rect 13282 27847 13502 27875
rect 13977 27847 14064 27875
rect 14530 27847 14750 27875
rect 13282 27801 13310 27847
rect 14722 27838 14750 27847
rect 16834 27847 17054 27875
rect 28450 27847 28574 27875
rect 16834 27838 16862 27847
rect 14722 27810 16862 27838
rect 4162 27773 4862 27801
rect 4162 27727 4190 27773
rect 34 27699 4190 27727
rect 4834 27727 4862 27773
rect 7522 27773 8414 27801
rect 12802 27773 13310 27801
rect 24994 27773 25598 27801
rect 7522 27727 7550 27773
rect 4834 27699 7550 27727
rect 8386 27727 8414 27773
rect 24994 27727 25022 27773
rect 8386 27699 11294 27727
rect 11266 27653 11294 27699
rect 12130 27699 12542 27727
rect 12130 27653 12158 27699
rect 4258 27625 4574 27653
rect 4642 27625 4766 27653
rect 7618 27625 7934 27653
rect 8002 27625 8318 27653
rect 11266 27625 12158 27653
rect 12514 27579 12542 27699
rect 13570 27699 18686 27727
rect 20962 27699 25022 27727
rect 25570 27727 25598 27773
rect 25570 27699 28670 27727
rect 28834 27699 29150 27727
rect 13570 27653 13598 27699
rect 13090 27625 13598 27653
rect 13785 27625 13872 27653
rect 16953 27625 17040 27653
rect 25090 27625 25502 27653
rect 26050 27625 26078 27699
rect 13090 27579 13118 27625
rect 1474 27551 3038 27579
rect 4377 27551 4464 27579
rect 5698 27551 6206 27579
rect 6370 27551 7824 27579
rect 12514 27551 13118 27579
rect 13762 27551 15696 27579
rect 17314 27551 17438 27579
rect 23266 27551 24734 27579
rect 26448 27551 26558 27579
rect 17314 27505 17342 27551
rect 4162 27477 4670 27505
rect 10018 27477 11102 27505
rect 16738 27477 17342 27505
rect 27106 27477 29726 27505
rect 10018 27431 10046 27477
rect 1954 27403 2846 27431
rect 3202 27403 3518 27431
rect 4258 27403 4958 27431
rect 9826 27403 10046 27431
rect 11074 27431 11102 27477
rect 24130 27440 26750 27468
rect 24130 27431 24158 27440
rect 11074 27403 11294 27431
rect 11458 27403 11870 27431
rect 13282 27403 13694 27431
rect 14722 27403 15230 27431
rect 23673 27403 23760 27431
rect 23938 27403 24158 27431
rect 26722 27431 26750 27440
rect 27106 27431 27134 27477
rect 26722 27403 27134 27431
rect 29698 27431 29726 27477
rect 29698 27403 29918 27431
rect 0 27257 32064 27355
rect 1570 27181 1982 27209
rect 6274 27181 6398 27209
rect 9634 27181 9854 27209
rect 6274 27061 6302 27181
rect 2434 27033 2544 27061
rect 4080 27033 6302 27061
rect 8002 27033 11678 27061
rect 11746 27033 14750 27061
rect 1282 26959 1406 26987
rect 1666 26959 2174 26987
rect 1666 26913 1694 26959
rect 1186 26885 1694 26913
rect 2146 26913 2174 26959
rect 2146 26885 2366 26913
rect 2722 26811 2750 26987
rect 7522 26959 7934 26987
rect 8025 26959 8112 26987
rect 9369 26959 9456 26987
rect 11746 26959 11774 27033
rect 11856 26959 11943 26987
rect 7906 26913 7934 26959
rect 12034 26913 12062 26987
rect 7906 26885 8702 26913
rect 9177 26885 9854 26913
rect 10882 26885 11582 26913
rect 11650 26885 12062 26913
rect 20889 26885 20976 26913
rect 21154 26885 21662 26913
rect 21826 26811 22334 26839
rect 21826 26802 21854 26811
rect 1954 26774 2558 26802
rect 1954 26765 1982 26774
rect 1762 26737 1982 26765
rect 2530 26765 2558 26774
rect 8482 26774 9182 26802
rect 8482 26765 8510 26774
rect 2530 26737 4670 26765
rect 5026 26737 5630 26765
rect 8290 26737 8510 26765
rect 9154 26765 9182 26774
rect 21058 26774 21854 26802
rect 21058 26765 21086 26774
rect 9154 26737 9374 26765
rect 20866 26737 21086 26765
rect 22306 26765 22334 26811
rect 22306 26737 22526 26765
rect 31234 26737 32030 26765
rect 0 26591 32064 26689
rect 13570 26515 13886 26543
rect 16546 26515 16766 26543
rect 20482 26515 20702 26543
rect 23746 26515 24446 26543
rect 29122 26515 29246 26543
rect 5506 26478 6014 26506
rect 5506 26469 5534 26478
rect 34 26441 254 26469
rect 226 26395 254 26441
rect 3682 26441 5534 26469
rect 5986 26469 6014 26478
rect 20482 26469 20510 26515
rect 5986 26441 10046 26469
rect 3682 26395 3710 26441
rect 10018 26395 10046 26441
rect 12034 26441 13790 26469
rect 12034 26395 12062 26441
rect 13762 26395 13790 26441
rect 14530 26441 16670 26469
rect 14530 26395 14558 26441
rect 226 26367 3710 26395
rect 4546 26367 4670 26395
rect 5602 26367 5918 26395
rect 8098 26367 8318 26395
rect 10018 26367 12062 26395
rect 13282 26367 13406 26395
rect 5602 26321 5630 26367
rect 3874 26293 4286 26321
rect 4354 26247 4382 26321
rect 4450 26293 5630 26321
rect 5890 26321 5918 26367
rect 5890 26293 6974 26321
rect 7138 26293 7934 26321
rect 8482 26293 8702 26321
rect 13570 26247 13598 26395
rect 13762 26367 14558 26395
rect 16642 26395 16670 26441
rect 18274 26441 18590 26469
rect 19810 26441 20510 26469
rect 18274 26395 18302 26441
rect 16642 26367 18302 26395
rect 19810 26321 19838 26441
rect 25378 26367 27422 26395
rect 28546 26367 31934 26395
rect 25378 26321 25406 26367
rect 14722 26293 14942 26321
rect 4354 26219 4574 26247
rect 4546 26210 4574 26219
rect 5314 26219 5534 26247
rect 7810 26219 8304 26247
rect 12226 26219 13598 26247
rect 14914 26247 14942 26293
rect 15874 26293 16094 26321
rect 16354 26293 16478 26321
rect 18466 26293 19838 26321
rect 19906 26293 20126 26321
rect 15874 26247 15902 26293
rect 14914 26219 15902 26247
rect 20098 26247 20126 26293
rect 20578 26293 22800 26321
rect 25186 26293 25406 26321
rect 27394 26321 27422 26367
rect 27394 26293 27600 26321
rect 20578 26247 20606 26293
rect 20098 26219 20606 26247
rect 22882 26219 23006 26247
rect 23097 26219 23184 26247
rect 24226 26219 26750 26247
rect 27609 26219 27696 26247
rect 27778 26219 27998 26247
rect 28953 26219 29040 26247
rect 5314 26210 5342 26219
rect 4546 26182 5342 26210
rect 22978 26173 23006 26219
rect 26722 26173 26750 26219
rect 27778 26173 27806 26219
rect 6274 26145 6974 26173
rect 22978 26145 23966 26173
rect 26722 26145 27806 26173
rect 3970 26071 4286 26099
rect 4930 26071 5726 26099
rect 6082 26071 6494 26099
rect 10233 26071 10320 26099
rect 16089 26071 16176 26099
rect 19353 26071 19440 26099
rect 0 25925 32064 26023
rect 6178 25849 7838 25877
rect 8098 25849 8318 25877
rect 9369 25849 9456 25877
rect 9634 25849 10718 25877
rect 16377 25849 16464 25877
rect 18658 25849 18878 25877
rect 18850 25803 18878 25849
rect 19714 25849 19934 25877
rect 21634 25849 21758 25877
rect 19714 25803 19742 25849
rect 18850 25775 19742 25803
rect 6850 25738 8222 25766
rect 6850 25729 6878 25738
rect 6658 25701 6878 25729
rect 8194 25729 8222 25738
rect 8194 25701 11294 25729
rect 11362 25701 13022 25729
rect 14818 25701 16670 25729
rect 20121 25701 20208 25729
rect 20386 25701 20510 25729
rect 21538 25701 23198 25729
rect 23650 25701 25392 25729
rect 729 25627 816 25655
rect 1186 25627 1406 25655
rect 1378 25618 1406 25627
rect 2530 25627 2750 25655
rect 6393 25627 8126 25655
rect 11362 25627 11390 25701
rect 11472 25627 11559 25655
rect 11664 25627 11751 25655
rect 14457 25627 14544 25655
rect 14841 25627 14928 25655
rect 18393 25627 18974 25655
rect 19426 25627 20112 25655
rect 25474 25627 25598 25655
rect 2530 25618 2558 25627
rect 1378 25590 2558 25618
rect 34 25553 638 25581
rect 610 25507 638 25553
rect 2818 25553 11294 25581
rect 2818 25507 2846 25553
rect 11266 25507 11294 25553
rect 11842 25553 18014 25581
rect 25186 25553 26462 25581
rect 11842 25507 11870 25553
rect 610 25479 2846 25507
rect 10809 25479 10896 25507
rect 11266 25479 11870 25507
rect 6754 25442 8222 25470
rect 6754 25433 6782 25442
rect 3033 25405 3120 25433
rect 6562 25405 6782 25433
rect 8194 25433 8222 25442
rect 8578 25442 10622 25470
rect 8578 25433 8606 25442
rect 8194 25405 8606 25433
rect 10594 25433 10622 25442
rect 14626 25442 15998 25470
rect 14626 25433 14654 25442
rect 10594 25405 11102 25433
rect 14434 25405 14654 25433
rect 15970 25433 15998 25442
rect 15970 25405 16286 25433
rect 27298 25405 27518 25433
rect 0 25259 32064 25357
rect 4066 25183 4286 25211
rect 14338 25183 14942 25211
rect 20098 25183 20414 25211
rect 20386 25137 20414 25183
rect 25090 25183 25694 25211
rect 26361 25183 26448 25211
rect 27778 25183 27998 25211
rect 22114 25146 24062 25174
rect 22114 25137 22142 25146
rect 4450 25109 4958 25137
rect 5794 25109 8318 25137
rect 20386 25109 22142 25137
rect 24034 25137 24062 25146
rect 25090 25137 25118 25183
rect 24034 25109 25118 25137
rect 25666 25137 25694 25183
rect 25666 25109 26270 25137
rect 3106 24961 4094 24989
rect 4066 24915 4094 24961
rect 4258 24961 4382 24989
rect 4450 24961 4478 25109
rect 5794 25063 5822 25109
rect 8290 25063 8318 25109
rect 4569 25035 5822 25063
rect 5913 25035 6000 25063
rect 6082 25035 6302 25063
rect 8098 25035 8222 25063
rect 8290 25035 8510 25063
rect 9346 25035 10238 25063
rect 10402 25035 11966 25063
rect 14361 25035 14448 25063
rect 15682 25035 16670 25063
rect 6082 24989 6110 25035
rect 4546 24961 4766 24989
rect 4258 24915 4286 24961
rect 1858 24887 2750 24915
rect 4066 24887 4286 24915
rect 4738 24915 4766 24961
rect 5602 24961 6110 24989
rect 5602 24915 5630 24961
rect 4738 24887 5630 24915
rect 6178 24915 6206 24989
rect 8313 24961 8400 24989
rect 9346 24915 9374 25035
rect 6178 24887 9374 24915
rect 10210 24915 10238 25035
rect 16642 24989 16670 25035
rect 22306 25035 23870 25063
rect 22306 24989 22334 25035
rect 10521 24961 10608 24989
rect 10704 24961 10791 24989
rect 12034 24961 12158 24989
rect 12240 24961 12327 24989
rect 12418 24915 12446 24989
rect 10210 24887 10526 24915
rect 10978 24887 12446 24915
rect 14242 24915 14270 24989
rect 16450 24961 16574 24989
rect 16642 24961 16766 24989
rect 21634 24961 22334 24989
rect 22402 24961 22526 24989
rect 23842 24915 23870 25035
rect 25282 25035 25502 25063
rect 25282 24915 25310 25035
rect 26242 24989 26270 25109
rect 27970 25063 27998 25183
rect 29986 25183 30206 25211
rect 29986 25137 30014 25183
rect 28738 25109 30014 25137
rect 31426 25109 31838 25137
rect 28738 25063 28766 25109
rect 31426 25063 31454 25109
rect 26352 25035 26439 25063
rect 27970 25035 28766 25063
rect 30370 25035 31454 25063
rect 30370 24989 30398 25035
rect 26242 24961 26558 24989
rect 30274 24961 30398 24989
rect 30466 24915 30494 24989
rect 30576 24961 30663 24989
rect 14242 24887 14366 24915
rect 19138 24887 20688 24915
rect 22224 24887 23678 24915
rect 23842 24887 25310 24915
rect 28930 24887 30110 24915
rect 30466 24887 30782 24915
rect 1858 24767 1886 24887
rect 1666 24739 1886 24767
rect 2722 24767 2750 24887
rect 9634 24776 11678 24804
rect 9634 24767 9662 24776
rect 2722 24739 2942 24767
rect 5794 24739 6014 24767
rect 8194 24739 8318 24767
rect 9442 24739 9662 24767
rect 11650 24767 11678 24776
rect 28930 24767 28958 24887
rect 11650 24739 11870 24767
rect 14050 24739 14174 24767
rect 16642 24739 16862 24767
rect 25858 24739 26078 24767
rect 28738 24739 28958 24767
rect 30082 24767 30110 24887
rect 30082 24739 30782 24767
rect 0 24593 32064 24691
rect 802 24517 1598 24545
rect 5794 24517 6014 24545
rect 6850 24517 7070 24545
rect 7042 24471 7070 24517
rect 7714 24517 8126 24545
rect 11074 24517 11582 24545
rect 14242 24517 14462 24545
rect 25762 24517 25886 24545
rect 7714 24471 7742 24517
rect 7042 24443 7742 24471
rect 7906 24443 8222 24471
rect 13282 24443 14558 24471
rect 18946 24443 19166 24471
rect 4546 24369 5630 24397
rect 8194 24383 8222 24443
rect 19138 24397 19166 24443
rect 19714 24443 21278 24471
rect 19714 24397 19742 24443
rect 21250 24397 21278 24443
rect 27202 24443 27614 24471
rect 27202 24397 27230 24443
rect 27586 24397 27614 24443
rect 28834 24443 29054 24471
rect 28834 24397 28862 24443
rect 19138 24369 19742 24397
rect 20313 24369 20400 24397
rect 21081 24369 21168 24397
rect 21250 24369 23486 24397
rect 25954 24369 26366 24397
rect 27010 24369 27230 24397
rect 27312 24369 27399 24397
rect 27586 24369 28862 24397
rect 4546 24323 4574 24369
rect 1378 24295 1694 24323
rect 4354 24295 4574 24323
rect 5602 24323 5630 24369
rect 5602 24295 6686 24323
rect 6873 24295 6960 24323
rect 7042 24295 8702 24323
rect 8674 24286 8702 24295
rect 9250 24295 9470 24323
rect 9250 24286 9278 24295
rect 8674 24258 9278 24286
rect 1209 24221 1296 24249
rect 1858 24221 2750 24249
rect 4162 24221 4286 24249
rect 4377 24221 4464 24249
rect 5602 24221 5726 24249
rect 1858 24101 1886 24221
rect 1666 24073 1886 24101
rect 2722 24101 2750 24221
rect 4258 24175 4286 24221
rect 5890 24175 5918 24249
rect 9538 24175 9566 24323
rect 10786 24295 12062 24323
rect 12921 24295 13008 24323
rect 14146 24295 14270 24323
rect 14338 24295 15518 24323
rect 19906 24295 20592 24323
rect 22521 24295 22608 24323
rect 10786 24249 10814 24295
rect 9922 24221 10142 24249
rect 10594 24221 10814 24249
rect 12034 24249 12062 24295
rect 14338 24249 14366 24295
rect 12034 24221 14366 24249
rect 22786 24175 22814 24249
rect 4258 24147 6686 24175
rect 8674 24147 9566 24175
rect 11650 24147 11774 24175
rect 21634 24147 22814 24175
rect 10498 24110 11486 24138
rect 10498 24101 10526 24110
rect 2722 24073 2942 24101
rect 4258 24073 4382 24101
rect 7618 24073 7934 24101
rect 10306 24073 10526 24101
rect 11458 24101 11486 24110
rect 11458 24073 11966 24101
rect 15609 24073 15696 24101
rect 20121 24073 20208 24101
rect 24322 24073 24734 24101
rect 0 23927 32064 24025
rect 1474 23851 1694 23879
rect 1666 23805 1694 23851
rect 2626 23851 2846 23879
rect 2914 23851 3038 23879
rect 5698 23851 5918 23879
rect 2626 23805 2654 23851
rect 5890 23842 5918 23851
rect 6658 23851 6878 23879
rect 7906 23851 8126 23879
rect 6658 23842 6686 23851
rect 5890 23814 6686 23842
rect 8098 23842 8126 23851
rect 9538 23851 9758 23879
rect 10114 23851 10334 23879
rect 12034 23851 12734 23879
rect 29890 23851 30206 23879
rect 8098 23814 8990 23842
rect 1666 23777 2654 23805
rect 8962 23805 8990 23814
rect 9538 23805 9566 23851
rect 8962 23777 9566 23805
rect 4162 23703 4382 23731
rect 4450 23703 5822 23731
rect 6274 23703 6686 23731
rect 6754 23703 6974 23731
rect 7042 23657 7070 23731
rect 8290 23703 8510 23731
rect 8697 23703 8784 23731
rect 13378 23703 14462 23731
rect 16450 23703 16670 23731
rect 16834 23703 16958 23731
rect 30178 23703 31934 23731
rect 13378 23657 13406 23703
rect 1282 23629 1598 23657
rect 1570 23583 1598 23629
rect 2722 23629 3134 23657
rect 3874 23629 4286 23657
rect 7042 23629 8414 23657
rect 8674 23629 9470 23657
rect 9538 23629 10142 23657
rect 10306 23629 11294 23657
rect 11554 23629 11678 23657
rect 12706 23629 13406 23657
rect 14434 23657 14462 23703
rect 14434 23629 14846 23657
rect 15682 23629 16766 23657
rect 30178 23629 30206 23703
rect 30393 23629 30480 23657
rect 2722 23583 2750 23629
rect 7042 23583 7070 23629
rect 9538 23583 9566 23629
rect 30562 23583 30590 23657
rect 1570 23555 2750 23583
rect 5794 23555 7070 23583
rect 9250 23555 9566 23583
rect 11074 23555 11390 23583
rect 7065 23481 7152 23509
rect 6274 23444 6878 23472
rect 6274 23435 6302 23444
rect 4450 23407 4766 23435
rect 6082 23407 6302 23435
rect 6850 23435 6878 23444
rect 6850 23407 7358 23435
rect 9826 23407 9950 23435
rect 11746 23407 11870 23435
rect 12994 23407 13310 23435
rect 13474 23407 13502 23569
rect 15129 23555 15216 23583
rect 29026 23555 30590 23583
rect 17122 23481 17630 23509
rect 17122 23435 17150 23481
rect 16930 23407 17150 23435
rect 17602 23435 17630 23481
rect 17602 23407 17822 23435
rect 30274 23407 30782 23435
rect 0 23261 32064 23359
rect 3874 23185 4478 23213
rect 4642 23185 4862 23213
rect 1186 23111 4382 23139
rect 4354 22991 4382 23111
rect 4450 23065 4478 23185
rect 4834 23176 4862 23185
rect 6754 23185 6974 23213
rect 13282 23185 13694 23213
rect 14242 23185 14462 23213
rect 4834 23148 6206 23176
rect 6178 23139 6206 23148
rect 6754 23139 6782 23185
rect 6178 23111 6782 23139
rect 14434 23139 14462 23185
rect 15010 23185 15230 23213
rect 15490 23185 15710 23213
rect 22521 23185 22608 23213
rect 15010 23139 15038 23185
rect 14434 23111 15038 23139
rect 19522 23111 23198 23139
rect 23170 23065 23198 23111
rect 23842 23111 25214 23139
rect 25378 23111 26366 23139
rect 27106 23111 28574 23139
rect 23842 23065 23870 23111
rect 4450 23037 6014 23065
rect 9058 23037 12734 23065
rect 17794 23037 17918 23065
rect 23170 23037 23870 23065
rect 2722 22963 3038 22991
rect 3321 22963 3408 22991
rect 4354 22963 4478 22991
rect 4546 22963 4670 22991
rect 5506 22963 5534 23037
rect 25762 23000 26270 23028
rect 25762 22991 25790 23000
rect 13872 22963 13959 22991
rect 14050 22963 14174 22991
rect 17433 22963 17520 22991
rect 18946 22963 19166 22991
rect 21442 22963 21662 22991
rect 21442 22917 21470 22963
rect 34 22889 2654 22917
rect 2626 22843 2654 22889
rect 3490 22889 13790 22917
rect 3490 22843 3518 22889
rect 13762 22880 13790 22889
rect 14242 22889 18878 22917
rect 20194 22889 20894 22917
rect 21058 22889 21470 22917
rect 21634 22917 21662 22963
rect 22594 22963 22814 22991
rect 24057 22963 24144 22991
rect 24226 22963 24350 22991
rect 22594 22917 22622 22963
rect 24418 22917 24446 22991
rect 24610 22963 24830 22991
rect 21634 22889 22622 22917
rect 22905 22889 22992 22917
rect 24034 22889 24446 22917
rect 24802 22917 24830 22963
rect 25570 22963 25790 22991
rect 26242 22991 26270 23000
rect 26242 22963 27518 22991
rect 27874 22963 28286 22991
rect 28368 22963 28455 22991
rect 25570 22917 25598 22963
rect 24802 22889 25598 22917
rect 26050 22889 26174 22917
rect 28642 22889 31454 22917
rect 14242 22880 14270 22889
rect 13762 22852 14270 22880
rect 28642 22843 28670 22889
rect 2626 22815 3518 22843
rect 4162 22815 4286 22843
rect 26722 22815 27710 22843
rect 27874 22815 28670 22843
rect 31426 22843 31454 22889
rect 31426 22815 31646 22843
rect 26722 22769 26750 22815
rect 5410 22741 5534 22769
rect 13666 22741 14366 22769
rect 21154 22741 21278 22769
rect 24034 22741 24350 22769
rect 25785 22741 25872 22769
rect 26530 22741 26750 22769
rect 27682 22769 27710 22815
rect 27682 22741 27998 22769
rect 0 22595 32064 22693
rect 2914 22519 3038 22547
rect 3394 22519 3614 22547
rect 5913 22519 6000 22547
rect 6201 22519 6288 22547
rect 7906 22519 8702 22547
rect 9058 22519 9278 22547
rect 19810 22519 20126 22547
rect 20098 22473 20126 22519
rect 22402 22519 22622 22547
rect 22882 22519 23006 22547
rect 25378 22519 25886 22547
rect 27394 22519 27614 22547
rect 22402 22510 22430 22519
rect 21058 22482 22430 22510
rect 27586 22510 27614 22519
rect 28450 22519 28670 22547
rect 28450 22510 28478 22519
rect 27586 22482 28478 22510
rect 21058 22473 21086 22482
rect 17026 22445 17534 22473
rect 20098 22445 21086 22473
rect 24034 22445 25310 22473
rect 17026 22399 17054 22445
rect 25282 22436 25310 22445
rect 26050 22445 27134 22473
rect 26050 22436 26078 22445
rect 25282 22408 26078 22436
rect 27106 22399 27134 22445
rect 5410 22371 5630 22399
rect 5721 22371 5808 22399
rect 5890 22371 6110 22399
rect 6082 22325 6110 22371
rect 6274 22371 7646 22399
rect 7906 22371 8894 22399
rect 9250 22371 9854 22399
rect 10594 22371 11294 22399
rect 11842 22371 12446 22399
rect 14626 22371 17054 22399
rect 21250 22371 22142 22399
rect 24322 22371 24446 22399
rect 27106 22371 29054 22399
rect 6274 22325 6302 22371
rect 3298 22297 3422 22325
rect 6082 22297 6302 22325
rect 7810 22251 7838 22325
rect 7906 22297 7934 22371
rect 10594 22251 10622 22371
rect 11266 22325 11294 22371
rect 11266 22297 11486 22325
rect 12034 22297 12638 22325
rect 17026 22297 17054 22371
rect 17122 22297 17438 22325
rect 21634 22297 21758 22325
rect 23001 22297 23088 22325
rect 23458 22297 24158 22325
rect 24130 22251 24158 22297
rect 25570 22297 25776 22325
rect 28546 22297 28670 22325
rect 25570 22251 25598 22297
rect 28930 22251 28958 22325
rect 29026 22297 29054 22371
rect 3586 22223 4382 22251
rect 7810 22223 8126 22251
rect 8194 22223 10622 22251
rect 12240 22223 15696 22251
rect 19138 22223 20400 22251
rect 24130 22223 25598 22251
rect 25762 22223 26078 22251
rect 26265 22223 26352 22251
rect 26914 22223 27326 22251
rect 27874 22223 28958 22251
rect 3586 22103 3614 22223
rect 3202 22075 3614 22103
rect 4354 22103 4382 22223
rect 5698 22149 5822 22177
rect 4354 22075 4574 22103
rect 10210 22075 10334 22103
rect 15129 22075 15216 22103
rect 29122 22075 29246 22103
rect 0 21929 32064 22027
rect 5602 21853 6110 21881
rect 6274 21853 6974 21881
rect 802 21816 2558 21844
rect 802 21807 830 21816
rect 34 21779 830 21807
rect 2530 21807 2558 21816
rect 6946 21807 6974 21853
rect 7714 21853 7934 21881
rect 8025 21853 8112 21881
rect 14073 21853 14160 21881
rect 14265 21853 14352 21881
rect 16642 21853 16862 21881
rect 17026 21853 17150 21881
rect 21561 21853 21648 21881
rect 27225 21853 27518 21881
rect 7714 21807 7742 21853
rect 25186 21816 26750 21844
rect 25186 21807 25214 21816
rect 2530 21779 3230 21807
rect 3298 21779 4478 21807
rect 6946 21779 7742 21807
rect 10402 21779 13982 21807
rect 3202 21659 3230 21779
rect 5794 21705 6782 21733
rect 8674 21705 9278 21733
rect 9442 21705 10238 21733
rect 1090 21631 1406 21659
rect 1378 21585 1406 21631
rect 2530 21631 2750 21659
rect 3202 21631 3518 21659
rect 2530 21585 2558 21631
rect 706 21557 1214 21585
rect 1378 21557 2558 21585
rect 3490 21585 3518 21631
rect 4162 21631 4766 21659
rect 5337 21631 5424 21659
rect 5986 21631 6302 21659
rect 6466 21631 6494 21705
rect 8674 21659 8702 21705
rect 7138 21631 7262 21659
rect 7344 21631 7431 21659
rect 8482 21631 8702 21659
rect 9250 21659 9278 21705
rect 9250 21631 10142 21659
rect 10233 21631 10320 21659
rect 10402 21631 10430 21779
rect 13954 21733 13982 21779
rect 14434 21779 16478 21807
rect 18850 21779 18974 21807
rect 23458 21779 25214 21807
rect 26722 21807 26750 21816
rect 27490 21807 27518 21853
rect 26722 21779 26942 21807
rect 27490 21779 28574 21807
rect 14434 21733 14462 21779
rect 13954 21705 14462 21733
rect 19426 21668 19934 21696
rect 19426 21659 19454 21668
rect 10498 21631 10910 21659
rect 11458 21631 11582 21659
rect 11746 21631 12062 21659
rect 12729 21631 12816 21659
rect 12994 21631 13118 21659
rect 16642 21631 16862 21659
rect 18466 21631 19454 21659
rect 19906 21659 19934 21668
rect 19906 21631 20126 21659
rect 20217 21631 20304 21659
rect 22306 21631 23198 21659
rect 23458 21631 23486 21779
rect 23554 21631 24062 21659
rect 25090 21631 25406 21659
rect 25488 21631 25575 21659
rect 26530 21631 26558 21719
rect 4162 21585 4190 21631
rect 4738 21585 4766 21631
rect 26914 21585 26942 21779
rect 28738 21705 31262 21733
rect 28738 21631 28766 21705
rect 28930 21585 28958 21659
rect 29040 21631 29127 21659
rect 3490 21557 4190 21585
rect 4354 21557 4478 21585
rect 4560 21557 4647 21585
rect 4738 21557 5246 21585
rect 5218 21548 5246 21557
rect 6562 21557 7070 21585
rect 7618 21557 8318 21585
rect 6562 21548 6590 21557
rect 5218 21520 6590 21548
rect 7618 21511 7646 21557
rect 7426 21483 7646 21511
rect 8290 21511 8318 21557
rect 12802 21557 18206 21585
rect 19545 21557 19632 21585
rect 20386 21557 21278 21585
rect 23746 21557 25022 21585
rect 12802 21548 12830 21557
rect 11554 21520 12830 21548
rect 11554 21511 11582 21520
rect 24994 21511 25022 21557
rect 25666 21557 26270 21585
rect 26914 21557 30686 21585
rect 25666 21511 25694 21557
rect 8290 21483 11582 21511
rect 12898 21483 13022 21511
rect 18370 21483 18782 21511
rect 23650 21483 24158 21511
rect 24994 21483 25694 21511
rect 23650 21437 23678 21483
rect 3202 21409 3326 21437
rect 6370 21409 6974 21437
rect 11650 21409 13982 21437
rect 23170 21409 23678 21437
rect 24130 21409 24158 21483
rect 29218 21409 29630 21437
rect 0 21263 32064 21361
rect 3106 21067 3134 21215
rect 5337 21187 5424 21215
rect 6946 21187 7358 21215
rect 11650 21187 11870 21215
rect 20290 21187 20510 21215
rect 20482 21178 20510 21187
rect 21346 21187 21566 21215
rect 22594 21187 22814 21215
rect 21346 21178 21374 21187
rect 20482 21150 21374 21178
rect 22786 21178 22814 21187
rect 23650 21187 24926 21215
rect 23650 21178 23678 21187
rect 22786 21150 23678 21178
rect 24898 21178 24926 21187
rect 26626 21187 29438 21215
rect 26626 21178 26654 21187
rect 24898 21150 26654 21178
rect 29410 21141 29438 21187
rect 30178 21187 30398 21215
rect 30178 21141 30206 21187
rect 3970 21113 5630 21141
rect 5602 21067 5630 21113
rect 20098 21067 20126 21141
rect 28834 21113 29246 21141
rect 29410 21113 30206 21141
rect 28834 21104 28862 21113
rect 23842 21076 24734 21104
rect 23842 21067 23870 21076
rect 1570 21039 3134 21067
rect 3202 21039 4094 21067
rect 4258 21039 4382 21067
rect 5602 21039 5726 21067
rect 7522 21039 8126 21067
rect 8290 21039 9758 21067
rect 11961 21039 12048 21067
rect 12921 21039 13008 21067
rect 13090 21039 13310 21067
rect 18105 21039 18192 21067
rect 20098 21039 21374 21067
rect 21442 21039 23870 21067
rect 24706 21067 24734 21076
rect 26818 21076 28862 21104
rect 26818 21067 26846 21076
rect 24706 21039 24926 21067
rect 7522 20993 7550 21039
rect 4546 20965 5342 20993
rect 6754 20965 6878 20993
rect 6960 20965 7047 20993
rect 7330 20965 7550 20993
rect 8098 20993 8126 21039
rect 8098 20965 8702 20993
rect 9561 20965 9648 20993
rect 10786 20965 11966 20993
rect 12898 20965 14558 20993
rect 14640 20965 14727 20993
rect 17506 20965 18014 20993
rect 4546 20919 4574 20965
rect 4258 20891 4574 20919
rect 5314 20919 5342 20965
rect 14530 20919 14558 20965
rect 21442 20919 21470 21039
rect 24898 20919 24926 21039
rect 25666 21039 26174 21067
rect 26338 21039 26846 21067
rect 29026 21039 29246 21067
rect 25666 20919 25694 21039
rect 26722 20965 27600 20993
rect 29218 20919 29246 21039
rect 30370 21039 30782 21067
rect 30370 20993 30398 21039
rect 30082 20965 30398 20993
rect 30585 20965 30672 20993
rect 30082 20919 30110 20965
rect 5314 20891 6302 20919
rect 7065 20891 7152 20919
rect 14530 20891 14750 20919
rect 19618 20891 21470 20919
rect 23074 20891 23294 20919
rect 23961 20891 24048 20919
rect 24130 20891 24638 20919
rect 24898 20891 25694 20919
rect 27609 20891 27696 20919
rect 27778 20891 27998 20919
rect 28930 20891 29054 20919
rect 29218 20891 30110 20919
rect 8194 20854 9278 20882
rect 8194 20845 8222 20854
rect 1570 20817 2942 20845
rect 6946 20817 8222 20845
rect 9250 20845 9278 20854
rect 27778 20845 27806 20891
rect 9250 20817 9470 20845
rect 26050 20817 27806 20845
rect 30754 20817 30782 21039
rect 30946 20817 31166 20845
rect 1570 20771 1598 20817
rect 1378 20743 1598 20771
rect 2914 20771 2942 20817
rect 4354 20780 5246 20808
rect 4354 20771 4382 20780
rect 2914 20743 3134 20771
rect 4162 20743 4382 20771
rect 5218 20771 5246 20780
rect 5218 20743 5438 20771
rect 5529 20743 5616 20771
rect 6489 20743 6576 20771
rect 8290 20743 8606 20771
rect 8985 20743 9072 20771
rect 9538 20743 10334 20771
rect 11458 20743 11774 20771
rect 12130 20743 13022 20771
rect 23001 20743 23088 20771
rect 25858 20743 25982 20771
rect 30274 20743 31934 20771
rect 0 20597 32064 20695
rect 1113 20521 1200 20549
rect 1497 20521 1584 20549
rect 4450 20521 4670 20549
rect 226 20447 1022 20475
rect 994 20438 1022 20447
rect 1666 20447 3518 20475
rect 1666 20438 1694 20447
rect 994 20410 1694 20438
rect 3490 20401 3518 20447
rect 3970 20447 4190 20475
rect 3970 20401 3998 20447
rect 3490 20373 3998 20401
rect 1305 20299 1392 20327
rect 1666 20299 3326 20327
rect 4450 20299 4478 20521
rect 4642 20475 4670 20521
rect 8098 20521 8318 20549
rect 8985 20521 9072 20549
rect 17410 20521 17534 20549
rect 20098 20521 20606 20549
rect 8098 20512 8126 20521
rect 5890 20484 8126 20512
rect 12034 20484 13982 20512
rect 5890 20475 5918 20484
rect 12034 20475 12062 20484
rect 4642 20447 5918 20475
rect 8770 20447 11582 20475
rect 11842 20447 12062 20475
rect 13954 20475 13982 20484
rect 13954 20447 14174 20475
rect 6082 20373 6590 20401
rect 8770 20387 8798 20447
rect 8962 20373 10046 20401
rect 10018 20364 10046 20373
rect 11266 20373 11486 20401
rect 11266 20364 11294 20373
rect 10018 20336 11294 20364
rect 11554 20327 11582 20447
rect 14146 20401 14174 20447
rect 12130 20373 12350 20401
rect 12418 20373 12528 20401
rect 14146 20373 18000 20401
rect 18480 20373 20510 20401
rect 12418 20327 12446 20373
rect 20482 20327 20510 20373
rect 4642 20299 6110 20327
rect 7522 20299 8606 20327
rect 8674 20299 9566 20327
rect 9730 20299 9854 20327
rect 11554 20299 12446 20327
rect 12633 20299 12720 20327
rect 20482 20299 20976 20327
rect 226 20225 1118 20253
rect 226 20179 254 20225
rect 34 20151 254 20179
rect 1090 20179 1118 20225
rect 5698 20225 5918 20253
rect 5698 20179 5726 20225
rect 1090 20151 3998 20179
rect 5602 20151 5726 20179
rect 4546 20077 4958 20105
rect 5986 20077 6014 20253
rect 6082 20225 6110 20299
rect 8674 20253 8702 20299
rect 6201 20225 6288 20253
rect 8386 20225 8702 20253
rect 9058 20225 9278 20253
rect 8386 20179 8414 20225
rect 9346 20179 9374 20253
rect 9561 20225 9648 20253
rect 9922 20225 10142 20253
rect 15202 20225 16574 20253
rect 16738 20225 16862 20253
rect 18178 20225 19358 20253
rect 19449 20225 19536 20253
rect 6658 20151 8414 20179
rect 8674 20151 9374 20179
rect 10114 20179 10142 20225
rect 10114 20151 14654 20179
rect 14818 20114 16382 20142
rect 14818 20105 14846 20114
rect 14146 20077 14846 20105
rect 16354 20105 16382 20114
rect 19330 20105 19358 20225
rect 19714 20151 20222 20179
rect 19714 20105 19742 20151
rect 16354 20077 16670 20105
rect 19330 20077 19742 20105
rect 20194 20105 20222 20151
rect 20578 20151 22142 20179
rect 20578 20105 20606 20151
rect 20194 20077 20606 20105
rect 22114 20105 22142 20151
rect 22306 20105 22334 20253
rect 22402 20225 22526 20253
rect 22114 20077 22334 20105
rect 0 19931 32064 20029
rect 7065 19855 7152 19883
rect 8770 19855 10526 19883
rect 27298 19855 27902 19883
rect 4354 19781 7262 19809
rect 3010 19707 3902 19735
rect 3010 19633 3038 19707
rect 4546 19670 5246 19698
rect 4546 19661 4574 19670
rect 4354 19633 4574 19661
rect 5218 19661 5246 19670
rect 5218 19633 5438 19661
rect 5529 19633 5616 19661
rect 5698 19633 5726 19781
rect 5817 19707 5904 19735
rect 6946 19707 7070 19735
rect 7138 19707 7358 19735
rect 7426 19707 8126 19735
rect 8770 19707 8798 19855
rect 12226 19781 16478 19809
rect 9154 19744 9758 19772
rect 9154 19735 9182 19744
rect 8962 19707 9182 19735
rect 9730 19735 9758 19744
rect 12226 19735 12254 19781
rect 9730 19707 9950 19735
rect 12226 19707 12350 19735
rect 7330 19587 7358 19707
rect 8194 19633 8894 19661
rect 8962 19633 8990 19707
rect 12226 19661 12254 19707
rect 16450 19661 16478 19781
rect 25090 19781 25598 19809
rect 25090 19735 25118 19781
rect 23074 19707 23582 19735
rect 23650 19707 23774 19735
rect 24802 19707 25118 19735
rect 25570 19735 25598 19781
rect 27874 19735 27902 19855
rect 30178 19855 30398 19883
rect 30178 19735 30206 19855
rect 25570 19707 25886 19735
rect 27874 19707 30206 19735
rect 30562 19707 31070 19735
rect 30562 19661 30590 19707
rect 8194 19587 8222 19633
rect 3010 19559 3134 19587
rect 4546 19559 6782 19587
rect 7330 19559 8222 19587
rect 9058 19513 9086 19661
rect 9346 19633 9854 19661
rect 10018 19633 10718 19661
rect 12034 19633 12254 19661
rect 12322 19633 14750 19661
rect 16450 19633 16958 19661
rect 17026 19633 17342 19661
rect 25186 19633 25502 19661
rect 30466 19633 30590 19661
rect 10690 19573 10718 19633
rect 12322 19513 12350 19633
rect 30658 19587 30686 19661
rect 30768 19633 30855 19661
rect 3874 19485 4382 19513
rect 9058 19485 10622 19513
rect 3874 19439 3902 19485
rect 4354 19476 4382 19485
rect 10594 19476 10622 19485
rect 12130 19485 12350 19513
rect 12418 19513 12446 19587
rect 17136 19559 18782 19587
rect 30658 19559 30974 19587
rect 12418 19485 12734 19513
rect 13858 19485 14078 19513
rect 12130 19476 12158 19485
rect 4354 19448 5534 19476
rect 10594 19448 12158 19476
rect 3106 19411 3326 19439
rect 3682 19411 3902 19439
rect 5506 19439 5534 19448
rect 5506 19411 5726 19439
rect 13401 19411 13488 19439
rect 13762 19411 14270 19439
rect 23938 19411 24254 19439
rect 30946 19411 31358 19439
rect 0 19265 32064 19363
rect 5794 19189 6014 19217
rect 5986 19143 6014 19189
rect 8866 19189 9278 19217
rect 5986 19115 7742 19143
rect 7714 19069 7742 19115
rect 8866 19069 8894 19189
rect 3225 19041 3312 19069
rect 4354 19041 5630 19069
rect 7714 19041 8894 19069
rect 9250 19069 9278 19189
rect 11266 19189 11870 19217
rect 12514 19189 12734 19217
rect 16354 19189 17054 19217
rect 22306 19189 22430 19217
rect 24322 19189 24542 19217
rect 11266 19069 11294 19189
rect 24514 19180 24542 19189
rect 27106 19189 27326 19217
rect 27106 19180 27134 19189
rect 24514 19152 27134 19180
rect 12034 19115 12350 19143
rect 9250 19041 11294 19069
rect 4354 18995 4382 19041
rect 2722 18967 4382 18995
rect 5602 18995 5630 19041
rect 12322 18995 12350 19115
rect 14722 19115 15806 19143
rect 14722 19069 14750 19115
rect 14338 19041 14750 19069
rect 15778 19069 15806 19115
rect 17698 19115 19358 19143
rect 17698 19069 17726 19115
rect 15778 19041 15998 19069
rect 16930 19041 17726 19069
rect 19330 19069 19358 19115
rect 19330 19041 19742 19069
rect 21744 19041 22142 19069
rect 24226 19041 24446 19069
rect 24418 18995 24446 19041
rect 24898 19041 25118 19069
rect 28066 19041 28190 19069
rect 28857 19041 28944 19069
rect 29337 19041 29424 19069
rect 24898 18995 24926 19041
rect 5602 18967 7550 18995
rect 2722 18893 2750 18967
rect 1186 18819 2558 18847
rect 1186 18773 1214 18819
rect 994 18745 1214 18773
rect 2530 18773 2558 18819
rect 2914 18819 3614 18847
rect 2914 18773 2942 18819
rect 2530 18745 2942 18773
rect 3586 18773 3614 18819
rect 4450 18819 7742 18847
rect 4450 18773 4478 18819
rect 3586 18745 3806 18773
rect 4258 18745 4478 18773
rect 7714 18773 7742 18819
rect 8098 18819 8894 18847
rect 8098 18773 8126 18819
rect 7714 18745 8126 18773
rect 8866 18773 8894 18819
rect 9058 18773 9086 18995
rect 11458 18967 12062 18995
rect 12144 18967 12231 18995
rect 12322 18967 12542 18995
rect 14818 18967 15902 18995
rect 16162 18967 16286 18995
rect 24418 18967 24926 18995
rect 25401 18967 25488 18995
rect 13378 18893 14174 18921
rect 17817 18893 17904 18921
rect 20194 18893 20318 18921
rect 20400 18893 20487 18921
rect 22306 18893 24062 18921
rect 13378 18847 13406 18893
rect 13186 18819 13406 18847
rect 14146 18847 14174 18893
rect 22306 18847 22334 18893
rect 14146 18819 20126 18847
rect 20098 18810 20126 18819
rect 20578 18819 22334 18847
rect 24034 18847 24062 18893
rect 27010 18893 27902 18921
rect 27010 18847 27038 18893
rect 27874 18884 27902 18893
rect 29698 18893 31838 18921
rect 27874 18856 28574 18884
rect 24034 18819 27038 18847
rect 28546 18847 28574 18856
rect 29698 18847 29726 18893
rect 28546 18819 29726 18847
rect 31810 18847 31838 18893
rect 31810 18819 32030 18847
rect 20578 18810 20606 18819
rect 20098 18782 20606 18810
rect 8866 18745 9086 18773
rect 17410 18745 17534 18773
rect 27874 18745 28478 18773
rect 0 18599 32064 18697
rect 3298 18523 4574 18551
rect 4546 18514 4574 18523
rect 5698 18523 6398 18551
rect 5698 18514 5726 18523
rect 4546 18486 5726 18514
rect 6370 18477 6398 18523
rect 7138 18523 7358 18551
rect 9538 18523 9758 18551
rect 10978 18523 11198 18551
rect 7138 18477 7166 18523
rect 9538 18514 9566 18523
rect 8482 18486 9566 18514
rect 4281 18449 4368 18477
rect 5890 18449 6014 18477
rect 6370 18449 7166 18477
rect 8002 18449 8126 18477
rect 4089 18375 4176 18403
rect 4450 18375 5822 18403
rect 994 18301 2942 18329
rect 3874 18301 4286 18329
rect 5890 18301 5918 18449
rect 7618 18375 7934 18403
rect 8482 18329 8510 18486
rect 8962 18375 9278 18403
rect 9465 18375 9552 18403
rect 9730 18375 9758 18523
rect 11170 18514 11198 18523
rect 12322 18523 12542 18551
rect 13282 18523 13502 18551
rect 12322 18514 12350 18523
rect 11170 18486 12350 18514
rect 13474 18477 13502 18523
rect 14050 18523 14846 18551
rect 14050 18477 14078 18523
rect 13474 18449 14078 18477
rect 14818 18403 14846 18523
rect 16066 18523 16286 18551
rect 17337 18523 17424 18551
rect 29410 18523 30206 18551
rect 16066 18403 16094 18523
rect 26050 18449 28574 18477
rect 28546 18403 28574 18449
rect 11170 18375 12062 18403
rect 14242 18375 14462 18403
rect 14553 18375 14640 18403
rect 14818 18375 16094 18403
rect 17904 18375 17991 18403
rect 22210 18375 25022 18403
rect 28377 18375 28464 18403
rect 28546 18375 28670 18403
rect 30274 18375 31550 18403
rect 22210 18329 22238 18375
rect 5986 18301 6206 18329
rect 7330 18301 7838 18329
rect 8002 18301 8510 18329
rect 8985 18301 9374 18329
rect 9442 18301 9662 18329
rect 9753 18301 9840 18329
rect 10018 18301 10526 18329
rect 16857 18301 16944 18329
rect 17218 18301 17534 18329
rect 21634 18301 22238 18329
rect 24994 18329 25022 18375
rect 25666 18338 26654 18366
rect 25666 18329 25694 18338
rect 24994 18301 25694 18329
rect 26626 18329 26654 18338
rect 26626 18301 27614 18329
rect 30274 18301 30302 18375
rect 4738 18227 5726 18255
rect 6466 18227 7166 18255
rect 8482 18227 8510 18301
rect 9346 18255 9374 18301
rect 10018 18255 10046 18301
rect 9346 18227 10046 18255
rect 10498 18255 10526 18301
rect 30466 18255 30494 18329
rect 30562 18301 30686 18329
rect 10498 18227 11486 18255
rect 17602 18227 17822 18255
rect 6466 18181 6494 18227
rect 6274 18153 6494 18181
rect 7138 18181 7166 18227
rect 17794 18181 17822 18227
rect 19330 18227 20126 18255
rect 19330 18181 19358 18227
rect 7138 18153 9086 18181
rect 17794 18153 19358 18181
rect 22210 18144 22238 18241
rect 22402 18227 24350 18255
rect 24802 18227 24926 18255
rect 24994 18144 25022 18241
rect 30466 18227 30974 18255
rect 22210 18116 25022 18144
rect 27778 18153 28670 18181
rect 27778 18107 27806 18153
rect 3106 18079 3326 18107
rect 9634 18079 10430 18107
rect 16953 18079 17040 18107
rect 19714 18079 19934 18107
rect 20194 18079 20510 18107
rect 26626 18079 27038 18107
rect 27298 18079 27806 18107
rect 28642 18107 28670 18153
rect 28642 18079 28862 18107
rect 30754 18079 31358 18107
rect 0 17933 32064 18031
rect 921 17857 1008 17885
rect 7330 17857 10622 17885
rect 11961 17857 12048 17885
rect 24322 17857 24638 17885
rect 24898 17857 25118 17885
rect 5986 17783 7358 17811
rect 7330 17774 7358 17783
rect 9922 17783 10142 17811
rect 9922 17774 9950 17783
rect 7330 17746 9950 17774
rect 3024 17709 3518 17737
rect 6178 17672 7166 17700
rect 6178 17663 6206 17672
rect 2722 17635 2846 17663
rect 3609 17635 3696 17663
rect 4066 17635 4382 17663
rect 4450 17635 4766 17663
rect 4857 17635 4944 17663
rect 5890 17589 5918 17663
rect 5986 17635 6206 17663
rect 7138 17663 7166 17672
rect 10594 17663 10622 17857
rect 25090 17811 25118 17857
rect 26050 17857 26270 17885
rect 29410 17857 29534 17885
rect 26050 17811 26078 17857
rect 27970 17820 29054 17848
rect 27970 17811 27998 17820
rect 16066 17783 16766 17811
rect 19330 17783 20414 17811
rect 25090 17783 26078 17811
rect 26530 17783 27422 17811
rect 27778 17783 27998 17811
rect 29026 17811 29054 17820
rect 29026 17783 31934 17811
rect 16066 17737 16094 17783
rect 15586 17709 16094 17737
rect 16738 17737 16766 17783
rect 16738 17709 16958 17737
rect 23746 17709 24446 17737
rect 27202 17709 27326 17737
rect 27394 17723 27422 17783
rect 7138 17635 10334 17663
rect 10402 17635 10526 17663
rect 10594 17635 10910 17663
rect 11746 17635 11966 17663
rect 12057 17635 12144 17663
rect 13282 17635 14174 17663
rect 15586 17635 15614 17709
rect 16162 17635 16766 17663
rect 16930 17635 16958 17709
rect 17506 17635 19838 17663
rect 19906 17635 20318 17663
rect 16162 17589 16190 17635
rect 24418 17589 24446 17709
rect 25378 17635 25886 17663
rect 27513 17635 27600 17663
rect 25378 17589 25406 17635
rect 3129 17561 3216 17589
rect 5122 17561 5726 17589
rect 5890 17561 6782 17589
rect 5122 17515 5150 17561
rect 4354 17487 5150 17515
rect 5698 17515 5726 17561
rect 6754 17515 6782 17561
rect 6946 17561 7070 17589
rect 10041 17561 10128 17589
rect 6946 17515 6974 17561
rect 7522 17524 8030 17552
rect 7522 17515 7550 17524
rect 5698 17487 6110 17515
rect 6585 17487 6672 17515
rect 6754 17487 6974 17515
rect 7330 17487 7550 17515
rect 8002 17515 8030 17524
rect 10594 17515 10622 17589
rect 10713 17561 10800 17589
rect 13977 17561 14064 17589
rect 14242 17561 14366 17589
rect 15417 17561 16190 17589
rect 16642 17561 17918 17589
rect 21634 17561 22142 17589
rect 22114 17515 22142 17561
rect 23362 17561 23582 17589
rect 23746 17561 23870 17589
rect 24153 17561 24240 17589
rect 24418 17561 25406 17589
rect 25858 17589 25886 17635
rect 25858 17561 26078 17589
rect 26242 17561 32030 17589
rect 23362 17515 23390 17561
rect 8002 17487 9662 17515
rect 10594 17487 12734 17515
rect 14530 17487 15038 17515
rect 6082 17441 6110 17487
rect 14530 17441 14558 17487
rect 6082 17413 7934 17441
rect 8674 17413 8894 17441
rect 14242 17413 14558 17441
rect 15010 17441 15038 17487
rect 19810 17487 20318 17515
rect 22114 17487 23390 17515
rect 17122 17450 18014 17478
rect 17122 17441 17150 17450
rect 15010 17413 15230 17441
rect 15394 17413 15710 17441
rect 16930 17413 17150 17441
rect 17986 17441 18014 17450
rect 19810 17441 19838 17487
rect 17986 17413 18206 17441
rect 18946 17413 19070 17441
rect 19618 17413 19838 17441
rect 20290 17441 20318 17487
rect 20290 17413 21086 17441
rect 21442 17413 21758 17441
rect 25474 17413 25790 17441
rect 0 17267 32064 17365
rect 3129 17191 3216 17219
rect 4162 17191 4574 17219
rect 6562 17191 7934 17219
rect 9177 17191 9264 17219
rect 10114 17191 10718 17219
rect 11577 17191 11664 17219
rect 12633 17191 12720 17219
rect 24153 17191 24240 17219
rect 25186 17191 25502 17219
rect 30946 17191 31070 17219
rect 4162 17182 4190 17191
rect 3298 17154 4190 17182
rect 3298 17145 3326 17154
rect 3010 17117 3326 17145
rect 4354 17117 5342 17145
rect 7257 17117 7344 17145
rect 8866 17117 9566 17145
rect 11266 17117 12062 17145
rect 12514 17117 12734 17145
rect 3490 17043 4478 17071
rect 4450 16997 4478 17043
rect 6274 17043 7070 17071
rect 6274 16997 6302 17043
rect 3225 16969 3518 16997
rect 3490 16960 3518 16969
rect 4162 16969 4382 16997
rect 4450 16969 4862 16997
rect 6201 16969 6302 16997
rect 4162 16960 4190 16969
rect 3490 16932 4190 16960
rect 6370 16923 6398 16997
rect 7234 16923 7262 17071
rect 11266 17043 11294 17117
rect 12706 17071 12734 17117
rect 13282 17117 14846 17145
rect 15106 17117 15518 17145
rect 13282 17071 13310 17117
rect 12706 17043 13310 17071
rect 8290 16969 8414 16997
rect 8482 16969 8606 16997
rect 11458 16923 11486 16997
rect 14818 16969 14846 17117
rect 15490 17071 15518 17117
rect 15778 17117 17150 17145
rect 15778 17071 15806 17117
rect 15129 17043 15216 17071
rect 15298 17043 15422 17071
rect 15490 17043 15806 17071
rect 17122 17071 17150 17117
rect 17890 17071 17918 17145
rect 17122 17043 18302 17071
rect 21058 17043 21278 17071
rect 21369 17043 21456 17071
rect 24418 17043 25022 17071
rect 15010 16969 15504 16997
rect 16944 16969 17054 16997
rect 17890 16969 18206 16997
rect 18274 16969 18302 17043
rect 24418 16997 24446 17043
rect 19618 16969 20414 16997
rect 23856 16969 24446 16997
rect 24994 16997 25022 17043
rect 26818 17043 28574 17071
rect 24994 16969 25584 16997
rect 26818 16983 26846 17043
rect 28258 16969 28478 16997
rect 28546 16983 28574 17043
rect 30658 16969 30974 16997
rect 418 16895 3038 16923
rect 4642 16895 5822 16923
rect 6370 16895 7262 16923
rect 10498 16895 12158 16923
rect 15010 16909 15038 16969
rect 17026 16923 17054 16969
rect 19618 16923 19646 16969
rect 17026 16895 18096 16923
rect 19440 16895 19646 16923
rect 418 16775 446 16895
rect 3010 16849 3038 16895
rect 3010 16821 4478 16849
rect 4450 16812 4478 16821
rect 6370 16812 6398 16895
rect 20386 16849 20414 16969
rect 28450 16923 28478 16969
rect 20482 16895 23006 16923
rect 23362 16895 23870 16923
rect 23961 16895 24048 16923
rect 24130 16895 25406 16923
rect 26434 16895 26558 16923
rect 26626 16895 26750 16923
rect 26914 16895 28382 16923
rect 28450 16895 28670 16923
rect 29698 16895 29918 16923
rect 23842 16849 23870 16895
rect 24130 16849 24158 16895
rect 8482 16821 9086 16849
rect 16066 16821 16862 16849
rect 20386 16821 20606 16849
rect 23842 16821 24158 16849
rect 26530 16849 26558 16895
rect 26914 16849 26942 16895
rect 26530 16821 26942 16849
rect 4450 16784 6398 16812
rect 11458 16784 12542 16812
rect 11458 16775 11486 16784
rect 226 16747 446 16775
rect 8025 16747 8112 16775
rect 9826 16747 10814 16775
rect 11266 16747 11486 16775
rect 12514 16775 12542 16784
rect 16066 16775 16094 16821
rect 12514 16747 12734 16775
rect 15874 16747 16094 16775
rect 16834 16775 16862 16821
rect 18850 16784 19934 16812
rect 18850 16775 18878 16784
rect 16834 16747 17438 16775
rect 18658 16747 18878 16775
rect 19906 16775 19934 16784
rect 19906 16747 20126 16775
rect 21346 16747 21662 16775
rect 28162 16747 28286 16775
rect 30850 16747 31070 16775
rect 0 16601 32064 16699
rect 802 16525 1022 16553
rect 994 16516 1022 16525
rect 2530 16525 2750 16553
rect 4834 16525 5054 16553
rect 2530 16516 2558 16525
rect 994 16488 2558 16516
rect 5026 16479 5054 16525
rect 8194 16525 8510 16553
rect 8985 16525 9072 16553
rect 10306 16525 10526 16553
rect 18178 16525 18302 16553
rect 20098 16525 20414 16553
rect 21826 16525 22334 16553
rect 8194 16516 8222 16525
rect 6178 16488 8222 16516
rect 6178 16479 6206 16488
rect 5026 16451 6206 16479
rect 22306 16479 22334 16525
rect 23554 16525 23774 16553
rect 24802 16525 25022 16553
rect 23554 16516 23582 16525
rect 22978 16488 23582 16516
rect 24994 16516 25022 16525
rect 25666 16525 25886 16553
rect 25666 16516 25694 16525
rect 24994 16488 25694 16516
rect 22978 16479 23006 16488
rect 22306 16451 23006 16479
rect 34 16331 62 16405
rect 2832 16377 4382 16405
rect 4354 16331 4382 16377
rect 7906 16331 7934 16391
rect 8025 16377 8112 16405
rect 8290 16377 10992 16405
rect 12633 16377 12720 16405
rect 13666 16377 14270 16405
rect 14626 16377 15326 16405
rect 21922 16377 22142 16405
rect 8290 16331 8318 16377
rect 13666 16331 13694 16377
rect 14626 16331 14654 16377
rect 34 16303 1214 16331
rect 1186 16294 1214 16303
rect 2242 16303 2654 16331
rect 4354 16303 4670 16331
rect 4738 16303 5150 16331
rect 2242 16294 2270 16303
rect 1186 16266 2270 16294
rect 2530 16229 3806 16257
rect 2530 16183 2558 16229
rect 3778 16220 3806 16229
rect 3778 16192 4286 16220
rect 34 16155 2558 16183
rect 4258 16183 4286 16192
rect 4738 16183 4766 16303
rect 5122 16257 5150 16303
rect 5602 16303 6302 16331
rect 5602 16257 5630 16303
rect 6274 16294 6302 16303
rect 7042 16303 7262 16331
rect 7522 16303 7742 16331
rect 7906 16303 8318 16331
rect 9369 16303 9456 16331
rect 12249 16303 12336 16331
rect 13378 16303 13694 16331
rect 14338 16303 14654 16331
rect 15298 16331 15326 16377
rect 15298 16303 15518 16331
rect 17049 16303 17136 16331
rect 18274 16303 18494 16331
rect 18585 16303 18672 16331
rect 19330 16303 20222 16331
rect 21273 16303 21360 16331
rect 7042 16294 7070 16303
rect 6274 16266 7070 16294
rect 13378 16257 13406 16303
rect 14338 16257 14366 16303
rect 21442 16257 21470 16331
rect 21561 16303 21648 16331
rect 5122 16229 5630 16257
rect 9250 16229 9566 16257
rect 10978 16229 13406 16257
rect 13474 16183 13502 16257
rect 13570 16229 14366 16257
rect 15682 16229 16382 16257
rect 17506 16229 17822 16257
rect 19906 16229 20126 16257
rect 20386 16229 21470 16257
rect 22114 16257 22142 16377
rect 23170 16377 23390 16405
rect 23842 16377 26366 16405
rect 23170 16331 23198 16377
rect 22786 16303 23198 16331
rect 22786 16257 22814 16303
rect 22114 16229 22814 16257
rect 23746 16257 23774 16331
rect 23842 16303 23870 16377
rect 26050 16303 26270 16331
rect 26338 16303 26366 16377
rect 26050 16294 26078 16303
rect 24898 16266 26078 16294
rect 24898 16257 24926 16266
rect 23746 16229 24926 16257
rect 26242 16257 26270 16303
rect 26242 16229 30878 16257
rect 15682 16220 15710 16229
rect 15202 16192 15710 16220
rect 15202 16183 15230 16192
rect 4258 16155 4766 16183
rect 5794 16155 8510 16183
rect 13474 16155 14078 16183
rect 14626 16155 15230 16183
rect 16354 16183 16382 16229
rect 16354 16155 17438 16183
rect 25090 16155 25694 16183
rect 25090 16146 25118 16155
rect 24226 16118 25118 16146
rect 24226 16109 24254 16118
rect 3321 16081 3408 16109
rect 9250 16081 9374 16109
rect 15298 16081 16286 16109
rect 18754 16081 18878 16109
rect 22978 16081 23486 16109
rect 24034 16081 24254 16109
rect 25666 16109 25694 16155
rect 25666 16081 25886 16109
rect 25954 16081 26462 16109
rect 26530 16081 26750 16109
rect 0 15935 32064 16033
rect 5410 15859 5822 15887
rect 9826 15859 9950 15887
rect 14050 15859 14270 15887
rect 2434 15665 2462 15739
rect 5410 15665 5438 15859
rect 5794 15739 5822 15859
rect 14242 15850 14270 15859
rect 15106 15859 15326 15887
rect 17721 15859 17808 15887
rect 18274 15859 20126 15887
rect 29890 15859 30014 15887
rect 15106 15850 15134 15859
rect 7330 15822 9758 15850
rect 14242 15822 15134 15850
rect 7330 15739 7358 15822
rect 9730 15813 9758 15822
rect 9730 15785 13118 15813
rect 15682 15785 16958 15813
rect 5794 15711 7358 15739
rect 7618 15711 9278 15739
rect 13282 15711 14942 15739
rect 13282 15665 13310 15711
rect 2434 15637 2654 15665
rect 3010 15637 3134 15665
rect 4738 15637 5438 15665
rect 5506 15637 5630 15665
rect 7522 15637 8030 15665
rect 11938 15637 12734 15665
rect 12921 15637 13310 15665
rect 14914 15665 14942 15711
rect 15682 15665 15710 15785
rect 16930 15739 16958 15785
rect 17218 15785 18494 15813
rect 26242 15785 28382 15813
rect 17218 15739 17246 15785
rect 18466 15776 18494 15785
rect 18466 15748 19742 15776
rect 19714 15739 19742 15748
rect 16930 15711 17246 15739
rect 17337 15711 17424 15739
rect 17506 15711 17630 15739
rect 17890 15711 18302 15739
rect 19714 15711 20030 15739
rect 14914 15637 15710 15665
rect 4738 15591 4766 15637
rect 11938 15591 11966 15637
rect 12706 15591 12734 15637
rect 4354 15563 4766 15591
rect 9360 15563 11966 15591
rect 12130 15563 12638 15591
rect 12706 15563 12816 15591
rect 14352 15563 15038 15591
rect 15010 15517 15038 15563
rect 15778 15517 15806 15651
rect 17314 15637 18014 15665
rect 18082 15637 18110 15711
rect 18274 15665 18302 15711
rect 20002 15665 20030 15711
rect 20482 15711 21374 15739
rect 28162 15711 28286 15739
rect 28354 15711 28382 15785
rect 29410 15711 30302 15739
rect 20482 15665 20510 15711
rect 16546 15563 16766 15591
rect 15010 15489 15806 15517
rect 16738 15517 16766 15563
rect 17314 15517 17342 15637
rect 18178 15591 18206 15665
rect 18274 15637 18686 15665
rect 19138 15637 19262 15665
rect 19344 15637 19431 15665
rect 20002 15637 20510 15665
rect 21346 15665 21374 15711
rect 21346 15637 21854 15665
rect 21922 15637 22238 15665
rect 30009 15637 30096 15665
rect 30274 15637 30302 15711
rect 30370 15637 30686 15665
rect 17506 15563 18206 15591
rect 19234 15591 19262 15637
rect 30370 15591 30398 15637
rect 19234 15563 20030 15591
rect 20578 15563 20688 15591
rect 16738 15489 17342 15517
rect 22018 15517 22046 15577
rect 26338 15563 30398 15591
rect 22018 15489 23006 15517
rect 12418 15452 14654 15480
rect 12418 15443 12446 15452
rect 6777 15415 6864 15443
rect 12226 15415 12446 15443
rect 14626 15443 14654 15452
rect 14626 15415 14846 15443
rect 18562 15415 18686 15443
rect 19161 15415 19248 15443
rect 28450 15415 28574 15443
rect 30562 15415 30974 15443
rect 0 15269 32064 15367
rect 3010 15193 3134 15221
rect 15609 15193 15696 15221
rect 25858 15193 26078 15221
rect 26050 15147 26078 15193
rect 31810 15193 32030 15221
rect 633 15119 720 15147
rect 34 15045 3614 15073
rect 13186 15059 13214 15147
rect 17698 15119 17918 15147
rect 17890 15073 17918 15119
rect 21346 15119 23870 15147
rect 26050 15119 27134 15147
rect 21346 15073 21374 15119
rect 27106 15073 27134 15119
rect 31810 15073 31838 15193
rect 17890 15045 21374 15073
rect 24706 15045 25310 15073
rect 27106 15045 31838 15073
rect 802 14999 830 15045
rect 3586 14999 3614 15045
rect 24706 14999 24734 15045
rect 706 14925 734 14999
rect 802 14971 1022 14999
rect 1666 14925 1694 14999
rect 2073 14971 2160 14999
rect 3586 14971 4094 14999
rect 12633 14971 12720 14999
rect 12802 14971 13118 14999
rect 15801 14971 15888 14999
rect 16258 14971 16478 14999
rect 22978 14971 23088 14999
rect 24528 14971 24734 14999
rect 25282 14999 25310 15045
rect 25282 14971 25488 14999
rect 12802 14925 12830 14971
rect 706 14897 1694 14925
rect 3129 14897 3216 14925
rect 3298 14897 3422 14925
rect 4354 14897 6110 14925
rect 7906 14897 12830 14925
rect 21538 14897 22910 14925
rect 3298 14851 3326 14897
rect 22882 14851 22910 14897
rect 24226 14897 24542 14925
rect 24610 14897 24734 14925
rect 25282 14897 25406 14925
rect 25474 14897 25598 14925
rect 24226 14851 24254 14897
rect 2626 14823 3326 14851
rect 4258 14823 4478 14851
rect 22882 14823 24254 14851
rect 24514 14851 24542 14897
rect 25474 14851 25502 14897
rect 24514 14823 27326 14851
rect 14146 14749 14942 14777
rect 16377 14749 16464 14777
rect 22306 14749 22622 14777
rect 27321 14749 27408 14777
rect 0 14603 32064 14701
rect 5529 14527 5616 14555
rect 6082 14527 8894 14555
rect 9538 14527 11006 14555
rect 12057 14527 12144 14555
rect 12706 14527 12926 14555
rect 5122 14453 6014 14481
rect 7714 14416 8414 14444
rect 7714 14407 7742 14416
rect 4258 14379 5342 14407
rect 5410 14379 5534 14407
rect 6777 14379 6864 14407
rect 6969 14379 7056 14407
rect 7426 14379 7742 14407
rect 8386 14407 8414 14416
rect 8386 14379 8606 14407
rect 7234 14305 8126 14333
rect 8866 14305 8894 14527
rect 12898 14481 12926 14527
rect 14146 14527 14366 14555
rect 18850 14527 19550 14555
rect 19810 14527 19934 14555
rect 21058 14527 21950 14555
rect 23458 14527 23678 14555
rect 14146 14481 14174 14527
rect 18850 14481 18878 14527
rect 12898 14453 14174 14481
rect 18178 14453 18878 14481
rect 10114 14416 10718 14444
rect 10114 14407 10142 14416
rect 9922 14379 10142 14407
rect 10690 14407 10718 14416
rect 10690 14379 10910 14407
rect 16258 14379 18110 14407
rect 10882 14333 10910 14379
rect 18178 14333 18206 14453
rect 9826 14305 10814 14333
rect 10882 14305 11006 14333
rect 11938 14305 12062 14333
rect 12921 14305 13008 14333
rect 13113 14305 13406 14333
rect 10882 14259 10910 14305
rect 13378 14259 13406 14305
rect 13954 14305 14558 14333
rect 14626 14305 14846 14333
rect 15682 14305 16190 14333
rect 13954 14259 13982 14305
rect 14626 14259 14654 14305
rect 34 14231 6302 14259
rect 7906 14231 8222 14259
rect 10594 14231 10910 14259
rect 11554 14231 13118 14259
rect 13378 14231 13982 14259
rect 14146 14231 14654 14259
rect 16162 14259 16190 14305
rect 17602 14305 17822 14333
rect 17890 14305 18206 14333
rect 19330 14333 19358 14481
rect 19330 14305 19454 14333
rect 19522 14305 19550 14527
rect 23650 14518 23678 14527
rect 24418 14527 24638 14555
rect 25378 14527 25598 14555
rect 29817 14527 29904 14555
rect 24418 14518 24446 14527
rect 23650 14490 24446 14518
rect 20098 14379 20894 14407
rect 21154 14379 21278 14407
rect 21826 14379 23294 14407
rect 23554 14379 25886 14407
rect 27586 14379 28478 14407
rect 25858 14333 25886 14379
rect 19618 14305 19742 14333
rect 20889 14305 20976 14333
rect 21346 14305 21758 14333
rect 22978 14305 23390 14333
rect 25474 14305 25790 14333
rect 25858 14305 25982 14333
rect 27682 14305 27998 14333
rect 17602 14259 17630 14305
rect 19618 14259 19646 14305
rect 16162 14231 17630 14259
rect 18754 14231 19646 14259
rect 26338 14231 27230 14259
rect 18754 14185 18782 14231
rect 18178 14157 18782 14185
rect 24514 14157 25982 14185
rect 24514 14111 24542 14157
rect 4546 14083 5438 14111
rect 5506 14083 6206 14111
rect 7234 14083 7358 14111
rect 8098 14083 8894 14111
rect 9561 14083 9648 14111
rect 11554 14083 12254 14111
rect 14722 14083 15326 14111
rect 17794 14083 18302 14111
rect 19042 14083 19262 14111
rect 21730 14083 21854 14111
rect 24322 14083 24542 14111
rect 25954 14111 25982 14157
rect 26338 14111 26366 14231
rect 25954 14083 26366 14111
rect 27202 14111 27230 14231
rect 27202 14083 27422 14111
rect 0 13937 32064 14035
rect 2073 13861 2160 13889
rect 6969 13861 7056 13889
rect 10233 13861 10320 13889
rect 11362 13861 13214 13889
rect 17721 13861 17808 13889
rect 21177 13861 21264 13889
rect 21826 13861 22046 13889
rect 22018 13852 22046 13861
rect 22978 13861 23198 13889
rect 26722 13861 26942 13889
rect 22978 13852 23006 13861
rect 22018 13824 23006 13852
rect 26914 13852 26942 13861
rect 31810 13861 32030 13889
rect 26914 13824 27806 13852
rect 27778 13815 27806 13824
rect 7906 13787 9470 13815
rect 11961 13787 12446 13815
rect 7906 13741 7934 13787
rect 1113 13713 1200 13741
rect 1378 13713 1694 13741
rect 1378 13667 1406 13713
rect 1666 13667 1694 13713
rect 3202 13713 3422 13741
rect 7714 13713 7934 13741
rect 9442 13741 9470 13787
rect 9442 13713 9662 13741
rect 3202 13667 3230 13713
rect 12418 13667 12446 13787
rect 15682 13787 17534 13815
rect 20674 13787 21566 13815
rect 27778 13787 29246 13815
rect 15682 13741 15710 13787
rect 29218 13741 29246 13787
rect 31810 13741 31838 13861
rect 13282 13713 15710 13741
rect 18658 13713 19166 13741
rect 20098 13713 20510 13741
rect 22114 13713 22430 13741
rect 23074 13713 24254 13741
rect 26530 13713 27614 13741
rect 29218 13713 31838 13741
rect 13282 13667 13310 13713
rect 18658 13667 18686 13713
rect 20482 13667 20510 13713
rect 22402 13667 22430 13713
rect 633 13639 720 13667
rect 1090 13639 1406 13667
rect 1474 13639 1598 13667
rect 1666 13639 1886 13667
rect 2626 13639 2846 13667
rect 3010 13639 3230 13667
rect 3298 13593 3326 13667
rect 3417 13639 3504 13667
rect 3586 13639 4478 13667
rect 5433 13639 5520 13667
rect 10329 13639 10416 13667
rect 11170 13639 11486 13667
rect 12418 13639 13310 13667
rect 16354 13639 16478 13667
rect 16546 13639 16766 13667
rect 3586 13593 3614 13639
rect 4450 13593 4478 13639
rect 16738 13593 16766 13639
rect 17602 13639 18686 13667
rect 19257 13639 19344 13667
rect 19906 13639 20414 13667
rect 20482 13639 21278 13667
rect 22210 13639 22334 13667
rect 22402 13639 23006 13667
rect 24418 13639 25790 13667
rect 25954 13639 26078 13667
rect 27586 13653 27614 13713
rect 17602 13593 17630 13639
rect 3202 13565 3614 13593
rect 4258 13565 4382 13593
rect 4450 13565 4574 13593
rect 4834 13565 5918 13593
rect 7906 13565 8030 13593
rect 10978 13565 11198 13593
rect 7906 13491 7934 13565
rect 11170 13519 11198 13565
rect 11362 13565 11966 13593
rect 12130 13565 12254 13593
rect 15874 13565 16190 13593
rect 16738 13565 17630 13593
rect 18009 13565 18096 13593
rect 19042 13565 19166 13593
rect 24322 13565 24542 13593
rect 25858 13565 27422 13593
rect 27490 13565 28286 13593
rect 11362 13519 11390 13565
rect 11170 13491 11390 13519
rect 19714 13491 21566 13519
rect 19714 13445 19742 13491
rect 3202 13417 3710 13445
rect 10690 13417 11102 13445
rect 16258 13417 16574 13445
rect 18082 13417 18878 13445
rect 19042 13417 19742 13445
rect 21538 13445 21566 13491
rect 28450 13491 29342 13519
rect 28450 13482 28478 13491
rect 26818 13454 28478 13482
rect 26818 13445 26846 13454
rect 21538 13417 21758 13445
rect 25858 13417 26270 13445
rect 26626 13417 26846 13445
rect 29314 13445 29342 13491
rect 29314 13417 29534 13445
rect 0 13271 32064 13369
rect 11458 13195 11678 13223
rect 11650 13149 11678 13195
rect 12706 13195 13214 13223
rect 12706 13149 12734 13195
rect 8098 13121 9374 13149
rect 11650 13121 12734 13149
rect 13186 13149 13214 13195
rect 13666 13195 13886 13223
rect 14530 13195 15134 13223
rect 15298 13195 15614 13223
rect 13666 13149 13694 13195
rect 13186 13121 13694 13149
rect 15586 13149 15614 13195
rect 16162 13195 16862 13223
rect 16162 13149 16190 13195
rect 15586 13121 16190 13149
rect 17890 13121 18782 13149
rect 19426 13121 20126 13149
rect 21538 13121 22142 13149
rect 8098 13075 8126 13121
rect 3586 13047 4094 13075
rect 5698 13047 5822 13075
rect 7833 13047 8126 13075
rect 3586 13001 3614 13047
rect 2434 12973 3614 13001
rect 4066 13001 4094 13047
rect 9346 13001 9374 13121
rect 9922 13047 10718 13075
rect 16377 13047 16464 13075
rect 18370 13047 18398 13121
rect 21538 13075 21566 13121
rect 18466 13047 18590 13075
rect 4066 12973 4862 13001
rect 9250 12927 9278 12987
rect 9346 12973 10334 13001
rect 12418 12973 12926 13001
rect 16473 12973 16560 13001
rect 12418 12927 12446 12973
rect 18658 12927 18686 13075
rect 18850 13047 18974 13075
rect 21346 13047 21566 13075
rect 22114 13075 22142 13121
rect 22114 13047 22334 13075
rect 22498 13047 23102 13075
rect 22498 13001 22526 13047
rect 21538 12973 22526 13001
rect 23074 13001 23102 13047
rect 23074 12973 23294 13001
rect 24610 12973 25214 13001
rect 24610 12927 24638 12973
rect 3682 12899 3998 12927
rect 5986 12899 6686 12927
rect 7138 12899 7646 12927
rect 9250 12899 10128 12927
rect 12130 12899 12446 12927
rect 13090 12899 13982 12927
rect 14146 12899 15038 12927
rect 15106 12899 18686 12927
rect 22128 12899 22238 12927
rect 22882 12899 23006 12927
rect 5986 12853 6014 12899
rect 5698 12825 6014 12853
rect 5698 12779 5726 12825
rect 4834 12751 5246 12779
rect 5506 12751 5726 12779
rect 6658 12779 6686 12899
rect 13090 12853 13118 12899
rect 10402 12825 10622 12853
rect 10594 12816 10622 12825
rect 11554 12825 12062 12853
rect 11554 12816 11582 12825
rect 10594 12788 11582 12816
rect 12034 12816 12062 12825
rect 12514 12825 13118 12853
rect 13954 12853 13982 12899
rect 22210 12853 22238 12899
rect 23074 12853 23102 12913
rect 24432 12899 24638 12927
rect 25186 12927 25214 12973
rect 25570 12973 26270 13001
rect 26553 12973 26640 13001
rect 27778 12973 28094 13001
rect 28162 12973 28286 13001
rect 25570 12927 25598 12973
rect 25186 12899 25598 12927
rect 26242 12927 26270 12973
rect 26242 12899 27984 12927
rect 31138 12899 31838 12927
rect 31138 12853 31166 12899
rect 13954 12825 14270 12853
rect 18274 12825 18494 12853
rect 22210 12825 23102 12853
rect 30946 12825 31166 12853
rect 31810 12853 31838 12899
rect 31810 12825 32030 12853
rect 12514 12816 12542 12825
rect 12034 12788 12542 12816
rect 28738 12788 29822 12816
rect 28738 12779 28766 12788
rect 6658 12751 6878 12779
rect 9657 12751 9744 12779
rect 14050 12751 14558 12779
rect 16738 12751 16958 12779
rect 24226 12751 25118 12779
rect 25666 12751 26366 12779
rect 28546 12751 28766 12779
rect 29794 12779 29822 12788
rect 29794 12751 30014 12779
rect 0 12605 32064 12703
rect 1474 12529 1790 12557
rect 5218 12529 5822 12557
rect 12034 12529 12350 12557
rect 12322 12520 12350 12529
rect 12898 12529 14366 12557
rect 15394 12529 16766 12557
rect 17506 12529 17726 12557
rect 12898 12520 12926 12529
rect 10210 12492 10718 12520
rect 12322 12492 12926 12520
rect 10210 12483 10238 12492
rect 1186 12455 1406 12483
rect 7330 12455 10238 12483
rect 10690 12483 10718 12492
rect 17698 12483 17726 12529
rect 18274 12529 18494 12557
rect 21154 12529 21374 12557
rect 22978 12529 23102 12557
rect 25785 12529 25872 12557
rect 28066 12529 28862 12557
rect 18274 12483 18302 12529
rect 10690 12455 11390 12483
rect 13090 12455 15134 12483
rect 15970 12455 17054 12483
rect 17698 12455 18302 12483
rect 1378 12446 1406 12455
rect 1378 12418 1982 12446
rect 130 12381 734 12409
rect 706 12335 734 12381
rect 1954 12335 1982 12418
rect 11650 12418 12158 12446
rect 11650 12409 11678 12418
rect 5122 12381 5726 12409
rect 10306 12381 11678 12409
rect 12130 12409 12158 12418
rect 12130 12381 13022 12409
rect 13282 12381 13598 12409
rect 5122 12335 5150 12381
rect 537 12307 624 12335
rect 706 12307 1790 12335
rect 1954 12307 2174 12335
rect 5026 12307 5150 12335
rect 5314 12307 5630 12335
rect 5314 12261 5342 12307
rect 3874 12233 4094 12261
rect 4546 12233 5342 12261
rect 5698 12261 5726 12381
rect 9657 12307 9744 12335
rect 10594 12307 11198 12335
rect 11746 12307 11870 12335
rect 12825 12307 12912 12335
rect 12994 12307 13022 12381
rect 13570 12335 13598 12381
rect 14242 12381 14462 12409
rect 20770 12381 21278 12409
rect 23938 12381 26846 12409
rect 28930 12381 29246 12409
rect 14242 12335 14270 12381
rect 13570 12307 14270 12335
rect 14818 12307 15710 12335
rect 16450 12307 16766 12335
rect 17794 12307 18110 12335
rect 18658 12307 19454 12335
rect 19522 12307 20702 12335
rect 20962 12307 22046 12335
rect 22114 12307 22910 12335
rect 25593 12307 25680 12335
rect 28258 12307 29054 12335
rect 18658 12261 18686 12307
rect 19522 12261 19550 12307
rect 5698 12233 6014 12261
rect 7042 12233 7646 12261
rect 8002 12233 9182 12261
rect 9442 12233 10430 12261
rect 11001 12233 11088 12261
rect 12802 12233 13406 12261
rect 18562 12233 18686 12261
rect 18754 12233 19550 12261
rect 22018 12261 22046 12307
rect 22018 12233 22814 12261
rect 22978 12233 23102 12261
rect 24226 12233 24350 12261
rect 25474 12233 25598 12261
rect 25858 12233 26270 12261
rect 27490 12233 28094 12261
rect 7042 12187 7070 12233
rect 6850 12159 7070 12187
rect 7618 12187 7646 12233
rect 7618 12159 7838 12187
rect 7810 12150 7838 12159
rect 9442 12159 9662 12187
rect 14050 12159 14558 12187
rect 9442 12150 9470 12159
rect 7810 12122 9470 12150
rect 12322 12122 13694 12150
rect 12322 12113 12350 12122
rect 2242 12085 2942 12113
rect 6178 12085 7166 12113
rect 12130 12085 12350 12113
rect 13666 12113 13694 12122
rect 14050 12113 14078 12159
rect 13666 12085 14078 12113
rect 14530 12113 14558 12159
rect 22210 12122 22814 12150
rect 22210 12113 22238 12122
rect 14530 12085 14750 12113
rect 17698 12085 18014 12113
rect 18754 12085 19070 12113
rect 19522 12085 19934 12113
rect 22018 12085 22238 12113
rect 22786 12113 22814 12122
rect 22978 12113 23006 12233
rect 27490 12187 27518 12233
rect 27298 12159 27518 12187
rect 28066 12187 28094 12233
rect 28066 12159 29438 12187
rect 22786 12085 23582 12113
rect 23746 12085 24254 12113
rect 0 11939 32064 12037
rect 7065 11863 7152 11891
rect 10329 11863 10416 11891
rect 10786 11863 11102 11891
rect 20985 11863 21072 11891
rect 23554 11863 23774 11891
rect 1378 11715 3902 11743
rect 5794 11715 6206 11743
rect 6969 11715 7056 11743
rect 7257 11715 7344 11743
rect 8985 11715 9072 11743
rect 130 11641 734 11669
rect 1113 11641 1200 11669
rect 4258 11641 5726 11669
rect 130 11493 158 11641
rect 5698 11595 5726 11641
rect 6274 11641 6590 11669
rect 6850 11641 7262 11669
rect 8793 11641 8880 11669
rect 10521 11641 10608 11669
rect 10786 11641 10814 11863
rect 11554 11789 13982 11817
rect 21922 11789 22142 11817
rect 13858 11669 13886 11743
rect 13954 11715 13982 11789
rect 23746 11743 23774 11863
rect 27682 11863 28094 11891
rect 27682 11743 27710 11863
rect 28066 11854 28094 11863
rect 28738 11863 28958 11891
rect 28738 11854 28766 11863
rect 28066 11826 28766 11854
rect 15394 11715 16574 11743
rect 16930 11715 17150 11743
rect 20674 11715 21086 11743
rect 21177 11715 21264 11743
rect 22018 11715 22526 11743
rect 23746 11715 27710 11743
rect 28162 11715 28574 11743
rect 15394 11669 15422 11715
rect 10896 11641 10983 11669
rect 12034 11641 12254 11669
rect 6274 11595 6302 11641
rect 12226 11595 12254 11641
rect 12994 11641 13406 11669
rect 13858 11641 14078 11669
rect 14242 11641 15422 11669
rect 16546 11669 16574 11715
rect 16546 11641 16766 11669
rect 22416 11641 22503 11669
rect 12994 11595 13022 11641
rect 537 11567 624 11595
rect 5698 11567 6302 11595
rect 8098 11567 8702 11595
rect 12226 11567 13022 11595
rect 13186 11567 13502 11595
rect 15490 11567 15600 11595
rect 18082 11567 21950 11595
rect 22320 11567 22407 11595
rect 20962 11456 21566 11484
rect 20962 11447 20990 11456
rect 1954 11419 2750 11447
rect 4642 11419 5054 11447
rect 8674 11419 9086 11447
rect 13186 11419 13598 11447
rect 14722 11419 14942 11447
rect 20313 11419 20400 11447
rect 20770 11419 20990 11447
rect 21538 11447 21566 11456
rect 21922 11456 22526 11484
rect 21922 11447 21950 11456
rect 21538 11419 21950 11447
rect 22498 11447 22526 11456
rect 22498 11419 23294 11447
rect 28066 11419 28286 11447
rect 0 11273 32064 11371
rect 1282 11197 1406 11225
rect 4761 11197 4848 11225
rect 8002 11197 8126 11225
rect 8793 11197 8880 11225
rect 9058 11151 9086 11225
rect 12825 11197 12912 11225
rect 13977 11197 14064 11225
rect 18658 11197 18878 11225
rect 18850 11151 18878 11197
rect 19330 11197 19550 11225
rect 20290 11197 20414 11225
rect 22402 11197 23198 11225
rect 23266 11197 24350 11225
rect 24610 11197 25022 11225
rect 19330 11151 19358 11197
rect 8194 11123 9086 11151
rect 11650 11123 16478 11151
rect 1570 11049 2366 11077
rect 1570 11003 1598 11049
rect 34 10975 1598 11003
rect 2338 11003 2366 11049
rect 11650 11003 11678 11123
rect 16450 11077 16478 11123
rect 17410 11123 17726 11151
rect 18850 11123 19358 11151
rect 17410 11077 17438 11123
rect 16450 11049 17438 11077
rect 17794 11049 18302 11077
rect 22498 11049 22718 11077
rect 2338 10975 8126 11003
rect 8098 10929 8126 10975
rect 9154 10975 11678 11003
rect 9154 10929 9182 10975
rect 13090 10929 13118 11003
rect 13762 10975 14366 11003
rect 14434 10975 15710 11003
rect 4281 10901 4368 10929
rect 8098 10901 9182 10929
rect 11746 10901 11870 10929
rect 11961 10901 12048 10929
rect 12994 10901 13118 10929
rect 13282 10901 13502 10929
rect 14626 10901 14750 10929
rect 13474 10855 13502 10901
rect 14722 10855 14750 10901
rect 15874 10855 15902 11003
rect 17794 10975 17822 11049
rect 22690 11003 22718 11049
rect 24034 11049 24542 11077
rect 24034 11003 24062 11049
rect 24514 11003 24542 11049
rect 25090 11049 26270 11077
rect 25090 11003 25118 11049
rect 19234 10975 19358 11003
rect 16066 10901 16286 10929
rect 17625 10901 17712 10929
rect 18082 10901 18206 10929
rect 19065 10901 19152 10929
rect 19234 10901 19262 10975
rect 20482 10929 20510 11003
rect 22690 10975 24062 11003
rect 24249 10975 24336 11003
rect 24514 10975 25118 11003
rect 19426 10901 20510 10929
rect 20674 10901 21086 10929
rect 26050 10901 26174 10929
rect 19426 10855 19454 10901
rect 1570 10827 2270 10855
rect 13378 10827 14558 10855
rect 14722 10827 15902 10855
rect 18466 10827 19454 10855
rect 1570 10781 1598 10827
rect 994 10753 1118 10781
rect 1378 10753 1598 10781
rect 2242 10781 2270 10827
rect 11938 10790 12542 10818
rect 11938 10781 11966 10790
rect 2242 10753 2462 10781
rect 3202 10753 3710 10781
rect 9849 10753 9936 10781
rect 11458 10753 11966 10781
rect 12514 10781 12542 10790
rect 12514 10753 12734 10781
rect 15970 10753 16286 10781
rect 18946 10753 19934 10781
rect 20482 10753 20606 10781
rect 23554 10753 24254 10781
rect 26361 10753 26448 10781
rect 0 10607 32064 10705
rect 1090 10531 1406 10559
rect 7042 10531 7166 10559
rect 9922 10531 10334 10559
rect 11170 10531 11582 10559
rect 12994 10531 13118 10559
rect 13186 10531 13310 10559
rect 15298 10531 16478 10559
rect 17026 10531 17726 10559
rect 25858 10531 26078 10559
rect 12034 10494 12830 10522
rect 12034 10485 12062 10494
rect 11842 10457 12062 10485
rect 12802 10485 12830 10494
rect 13090 10485 13118 10531
rect 13762 10494 14366 10522
rect 13762 10485 13790 10494
rect 12802 10457 13022 10485
rect 13090 10457 13790 10485
rect 14338 10485 14366 10494
rect 14338 10457 15230 10485
rect 11842 10411 11870 10457
rect 12994 10411 13022 10457
rect 15202 10448 15230 10457
rect 16066 10457 17150 10485
rect 18754 10457 19550 10485
rect 16066 10448 16094 10457
rect 15202 10420 16094 10448
rect 18754 10411 18782 10457
rect 19522 10411 19550 10457
rect 21442 10457 21662 10485
rect 26242 10457 26654 10485
rect 21442 10411 21470 10457
rect 26626 10411 26654 10457
rect 27202 10457 29822 10485
rect 31330 10457 32030 10485
rect 27202 10411 27230 10457
rect 6850 10383 7262 10411
rect 8098 10383 8702 10411
rect 8866 10383 9758 10411
rect 1113 10309 1200 10337
rect 1474 10309 1694 10337
rect 2434 10309 4574 10337
rect 4761 10309 4848 10337
rect 5122 10309 5246 10337
rect 7042 10309 7166 10337
rect 7234 10309 7262 10383
rect 8866 10337 8894 10383
rect 8194 10309 8894 10337
rect 9730 10337 9758 10383
rect 10786 10383 11870 10411
rect 12034 10383 12926 10411
rect 12994 10383 13214 10411
rect 10786 10337 10814 10383
rect 12034 10337 12062 10383
rect 13186 10374 13214 10383
rect 13858 10383 14270 10411
rect 16258 10383 17054 10411
rect 17986 10383 18782 10411
rect 19257 10383 19344 10411
rect 19522 10383 21470 10411
rect 23074 10383 23774 10411
rect 24130 10383 24254 10411
rect 26626 10383 27230 10411
rect 13858 10374 13886 10383
rect 13186 10346 13886 10374
rect 17986 10337 18014 10383
rect 9730 10309 10814 10337
rect 10882 10309 11006 10337
rect 11746 10309 12062 10337
rect 12994 10263 13022 10337
rect 994 10235 2366 10263
rect 2338 10226 2366 10235
rect 3010 10235 3230 10263
rect 3010 10226 3038 10235
rect 2338 10198 3038 10226
rect 9634 10189 9662 10249
rect 12034 10235 13022 10263
rect 13858 10235 13982 10263
rect 14050 10189 14078 10323
rect 17410 10309 18014 10337
rect 18873 10309 18960 10337
rect 19042 10309 19262 10337
rect 21922 10263 21950 10337
rect 23746 10309 23774 10383
rect 23961 10309 24048 10337
rect 27394 10309 27998 10337
rect 21730 10235 21950 10263
rect 22114 10235 25982 10263
rect 27586 10235 27710 10263
rect 18082 10198 18974 10226
rect 18082 10189 18110 10198
rect 9634 10161 11966 10189
rect 11938 10152 11966 10161
rect 13090 10161 14078 10189
rect 14530 10161 18110 10189
rect 18946 10189 18974 10198
rect 18946 10161 19166 10189
rect 23554 10161 23774 10189
rect 13090 10152 13118 10161
rect 11938 10124 13118 10152
rect 23554 10115 23582 10161
rect 2434 10087 3134 10115
rect 5890 10087 6398 10115
rect 10402 10087 10622 10115
rect 11673 10087 11760 10115
rect 17314 10087 17534 10115
rect 18178 10087 18878 10115
rect 22018 10087 22334 10115
rect 23266 10087 23582 10115
rect 23650 10087 23870 10115
rect 0 9941 32064 10039
rect 2146 9865 2366 9893
rect 2338 9856 2366 9865
rect 3298 9865 3902 9893
rect 12514 9865 12734 9893
rect 3298 9856 3326 9865
rect 2338 9828 3326 9856
rect 12706 9856 12734 9865
rect 17986 9865 18206 9893
rect 19330 9865 19742 9893
rect 17986 9856 18014 9865
rect 12706 9828 15806 9856
rect 15778 9819 15806 9828
rect 16930 9828 18014 9856
rect 19714 9856 19742 9865
rect 20674 9865 20894 9893
rect 23458 9865 23870 9893
rect 27682 9865 27806 9893
rect 20674 9856 20702 9865
rect 19714 9828 20702 9856
rect 16930 9819 16958 9828
rect 3490 9754 4094 9782
rect 3490 9745 3518 9754
rect 2722 9717 3518 9745
rect 4066 9745 4094 9754
rect 4066 9717 4958 9745
rect 7426 9717 7920 9745
rect 8386 9731 8414 9819
rect 15778 9791 16958 9819
rect 18274 9791 19550 9819
rect 27106 9791 27902 9819
rect 22978 9754 23582 9782
rect 22978 9745 23006 9754
rect 11554 9717 12734 9745
rect 1378 9643 1502 9671
rect 1762 9643 2462 9671
rect 1762 9569 1790 9643
rect 2530 9597 2558 9671
rect 3705 9643 3792 9671
rect 3970 9597 3998 9671
rect 7426 9657 7454 9717
rect 8098 9643 8222 9671
rect 9442 9643 11390 9671
rect 11472 9643 11559 9671
rect 11650 9643 11774 9671
rect 11362 9597 11390 9643
rect 1858 9569 1982 9597
rect 2050 9569 2558 9597
rect 3490 9569 3998 9597
rect 7257 9569 7344 9597
rect 7545 9569 7632 9597
rect 7714 9569 8030 9597
rect 11362 9569 11582 9597
rect 12706 9569 12734 9717
rect 17122 9717 18206 9745
rect 17122 9671 17150 9717
rect 13090 9643 15806 9671
rect 15778 9597 15806 9643
rect 16642 9643 17150 9671
rect 18178 9643 18206 9717
rect 18946 9717 21758 9745
rect 22498 9717 23006 9745
rect 23554 9745 23582 9754
rect 23554 9717 23774 9745
rect 27106 9731 27134 9791
rect 18274 9643 18398 9671
rect 16642 9597 16670 9643
rect 18946 9597 18974 9717
rect 19234 9643 19358 9671
rect 19449 9643 19536 9671
rect 12802 9569 12926 9597
rect 13008 9569 13095 9597
rect 15778 9569 16670 9597
rect 17314 9569 18974 9597
rect 5698 9495 6686 9523
rect 5698 9449 5726 9495
rect 1401 9421 1488 9449
rect 1666 9421 2270 9449
rect 3298 9421 4190 9449
rect 5506 9421 5726 9449
rect 6658 9449 6686 9495
rect 9250 9495 9758 9523
rect 11554 9495 11582 9569
rect 20464 9560 20528 9683
rect 21922 9643 22622 9671
rect 20578 9569 20702 9597
rect 21922 9569 21950 9643
rect 22594 9597 22622 9643
rect 23074 9643 23294 9671
rect 23746 9643 23774 9717
rect 29026 9717 29246 9745
rect 29026 9671 29054 9717
rect 26914 9643 27422 9671
rect 27970 9643 29054 9671
rect 29410 9643 29534 9671
rect 23074 9597 23102 9643
rect 22018 9523 22046 9597
rect 22137 9569 22224 9597
rect 22320 9569 22407 9597
rect 22594 9569 23102 9597
rect 23650 9569 23870 9597
rect 25378 9569 27326 9597
rect 27705 9569 27792 9597
rect 28066 9569 28286 9597
rect 11938 9495 12542 9523
rect 9250 9449 9278 9495
rect 6658 9421 6878 9449
rect 9058 9421 9278 9449
rect 9730 9449 9758 9495
rect 11938 9449 11966 9495
rect 12514 9486 12542 9495
rect 13282 9495 15422 9523
rect 18946 9495 22046 9523
rect 13282 9486 13310 9495
rect 12514 9458 13310 9486
rect 9730 9421 9950 9449
rect 10594 9421 11966 9449
rect 15394 9449 15422 9495
rect 17026 9458 17822 9486
rect 17026 9449 17054 9458
rect 15394 9421 15614 9449
rect 16834 9421 17054 9449
rect 17794 9449 17822 9458
rect 17794 9421 18014 9449
rect 20098 9421 20222 9449
rect 20290 9421 20414 9449
rect 23074 9421 23678 9449
rect 25017 9421 25104 9449
rect 0 9275 32064 9373
rect 1090 9199 1886 9227
rect 1977 9199 2064 9227
rect 2338 9199 3326 9227
rect 4546 9199 4766 9227
rect 5026 9199 5150 9227
rect 5794 9199 6206 9227
rect 7426 9199 7646 9227
rect 8002 9199 8126 9227
rect 11170 9199 11486 9227
rect 4738 9153 4766 9199
rect 11458 9190 11486 9199
rect 13666 9199 13886 9227
rect 13954 9199 14174 9227
rect 18082 9199 18302 9227
rect 19234 9199 19454 9227
rect 11458 9162 12350 9190
rect 12322 9153 12350 9162
rect 13666 9153 13694 9199
rect 14914 9162 15422 9190
rect 14914 9153 14942 9162
rect 2722 9125 3998 9153
rect 1186 9088 1790 9116
rect 1186 9079 1214 9088
rect 802 9051 1214 9079
rect 1762 9079 1790 9088
rect 1762 9051 2366 9079
rect 802 9005 830 9051
rect 2338 9005 2366 9051
rect 2722 9005 2750 9125
rect 4450 9079 4478 9153
rect 4738 9125 5726 9153
rect 5698 9116 5726 9125
rect 6274 9125 6494 9153
rect 6274 9116 6302 9125
rect 5698 9088 6302 9116
rect 3010 9051 3326 9079
rect 4450 9051 4958 9079
rect 3010 9005 3038 9051
rect 3298 9005 3326 9051
rect 130 8977 830 9005
rect 898 8977 1502 9005
rect 2338 8977 2750 9005
rect 2818 8977 3038 9005
rect 3106 8977 3230 9005
rect 3298 8977 3614 9005
rect 4089 8977 4176 9005
rect 4258 8977 4478 9005
rect 4560 8977 4647 9005
rect 4450 8931 4478 8977
rect 4738 8931 4766 9005
rect 4930 8977 4958 9051
rect 5986 8977 6206 9005
rect 6562 8977 6686 9005
rect 6850 8977 6974 9005
rect 7042 8977 7070 9153
rect 10498 9125 11294 9153
rect 12322 9125 13694 9153
rect 14146 9125 14942 9153
rect 15394 9153 15422 9162
rect 16834 9162 17438 9190
rect 16834 9153 16862 9162
rect 15394 9125 16862 9153
rect 17410 9153 17438 9162
rect 19426 9153 19454 9199
rect 19906 9199 20414 9227
rect 21058 9199 22430 9227
rect 19906 9153 19934 9199
rect 17410 9125 18206 9153
rect 19426 9125 19934 9153
rect 11266 9079 11294 9125
rect 8482 9051 9182 9079
rect 7161 8977 7248 9005
rect 5986 8931 6014 8977
rect 2928 8903 3015 8931
rect 4450 8903 4670 8931
rect 4738 8903 6014 8931
rect 1570 8829 2750 8857
rect 1570 8783 1598 8829
rect 2722 8820 2750 8829
rect 3874 8829 4862 8857
rect 2722 8792 3422 8820
rect 1378 8755 1598 8783
rect 3394 8783 3422 8792
rect 3874 8783 3902 8829
rect 5026 8783 5054 8903
rect 8290 8857 8318 9005
rect 8482 8977 8510 9051
rect 9346 9005 9374 9079
rect 10521 9051 10608 9079
rect 11266 9051 12158 9079
rect 14146 9005 14174 9125
rect 15010 9051 15326 9079
rect 16930 9051 17342 9079
rect 17986 9051 18110 9079
rect 19161 9051 19248 9079
rect 20386 9051 20414 9199
rect 22402 9153 22430 9199
rect 24610 9199 25118 9227
rect 25305 9199 25392 9227
rect 24610 9190 24638 9199
rect 23266 9162 24638 9190
rect 23266 9153 23294 9162
rect 20496 9125 20583 9153
rect 22402 9125 23294 9153
rect 26242 9079 26270 9153
rect 21730 9051 22142 9079
rect 15010 9005 15038 9051
rect 15298 9005 15326 9051
rect 21730 9005 21758 9051
rect 8578 8977 10142 9005
rect 10233 8977 10320 9005
rect 10402 8931 10430 9005
rect 10978 8977 11390 9005
rect 11481 8977 11568 9005
rect 11650 8977 14174 9005
rect 14242 8977 15038 9005
rect 15129 8977 15216 9005
rect 15298 8977 15518 9005
rect 15586 8977 16670 9005
rect 16738 8977 17246 9005
rect 18393 8977 18480 9005
rect 20674 8977 21758 9005
rect 17218 8931 17246 8977
rect 21826 8931 21854 9005
rect 22114 8977 22142 9051
rect 23554 9051 24158 9079
rect 25666 9051 26750 9079
rect 23554 9005 23582 9051
rect 23458 8977 23582 9005
rect 23664 8977 23751 9005
rect 24226 8977 25214 9005
rect 28258 8977 28670 9005
rect 28834 8977 28958 9005
rect 9634 8903 10910 8931
rect 11746 8903 11966 8931
rect 17218 8903 20318 8931
rect 21826 8903 23102 8931
rect 24226 8903 24254 8977
rect 25474 8903 26846 8931
rect 27010 8903 27614 8931
rect 10882 8857 10910 8903
rect 13858 8866 15422 8894
rect 13858 8857 13886 8866
rect 8290 8829 9278 8857
rect 10882 8829 13886 8857
rect 15394 8857 15422 8866
rect 27010 8857 27038 8903
rect 15394 8829 16382 8857
rect 26626 8829 27038 8857
rect 27586 8857 27614 8903
rect 27586 8829 28670 8857
rect 26626 8820 26654 8829
rect 25186 8792 26654 8820
rect 25186 8783 25214 8792
rect 3394 8755 3902 8783
rect 3970 8755 5054 8783
rect 13954 8755 15326 8783
rect 16450 8755 16862 8783
rect 18082 8755 18398 8783
rect 19449 8755 19536 8783
rect 21561 8755 21648 8783
rect 23481 8755 23568 8783
rect 24706 8755 25214 8783
rect 26722 8755 27038 8783
rect 0 8609 32064 8707
rect 1186 8533 1406 8561
rect 1378 8524 1406 8533
rect 2146 8533 2558 8561
rect 3778 8533 4670 8561
rect 6658 8533 6782 8561
rect 12729 8533 12816 8561
rect 13113 8533 13200 8561
rect 15129 8533 15216 8561
rect 16354 8533 16862 8561
rect 17506 8533 17918 8561
rect 19426 8533 19550 8561
rect 20674 8533 20894 8561
rect 21657 8533 21744 8561
rect 21922 8533 22142 8561
rect 22306 8533 23294 8561
rect 24610 8533 24734 8561
rect 25666 8533 25790 8561
rect 29602 8533 29822 8561
rect 2146 8524 2174 8533
rect 1378 8496 2174 8524
rect 2338 8459 3614 8487
rect 3586 8413 3614 8459
rect 4162 8459 4382 8487
rect 8866 8459 9278 8487
rect 4162 8413 4190 8459
rect 1762 8385 2846 8413
rect 3586 8385 4190 8413
rect 2818 8339 2846 8385
rect 2073 8311 2160 8339
rect 2338 8311 2750 8339
rect 2818 8311 3422 8339
rect 4354 8311 4478 8339
rect 4546 8311 5534 8339
rect 6946 8311 7742 8339
rect 8194 8311 8798 8339
rect 8866 8265 8894 8459
rect 9250 8413 9278 8459
rect 10114 8459 10334 8487
rect 12130 8459 13118 8487
rect 18466 8459 20126 8487
rect 22882 8459 24254 8487
rect 10114 8413 10142 8459
rect 22882 8413 22910 8459
rect 29794 8413 29822 8533
rect 31618 8533 31838 8561
rect 31618 8413 31646 8533
rect 9250 8385 10142 8413
rect 15394 8385 16766 8413
rect 15394 8339 15422 8385
rect 8985 8311 9072 8339
rect 12130 8311 12350 8339
rect 1090 8237 1502 8265
rect 2434 8191 2462 8265
rect 2553 8237 2640 8265
rect 5122 8237 6398 8265
rect 6466 8237 6590 8265
rect 8098 8237 8894 8265
rect 12322 8265 12350 8311
rect 12802 8311 13022 8339
rect 15010 8311 15422 8339
rect 16738 8339 16766 8385
rect 20482 8339 20510 8413
rect 21922 8385 22910 8413
rect 23362 8385 23486 8413
rect 25954 8385 28382 8413
rect 29794 8385 31646 8413
rect 21922 8339 21950 8385
rect 16738 8311 18110 8339
rect 18274 8311 18974 8339
rect 19426 8311 19550 8339
rect 20386 8311 20510 8339
rect 12802 8265 12830 8311
rect 12322 8237 12830 8265
rect 13305 8237 13392 8265
rect 15010 8237 15038 8311
rect 18274 8265 18302 8311
rect 15120 8237 15207 8265
rect 15298 8237 15422 8265
rect 16185 8237 16272 8265
rect 16354 8191 16382 8265
rect 16450 8237 16574 8265
rect 1570 8163 2462 8191
rect 14338 8163 16382 8191
rect 16642 8117 16670 8265
rect 17602 8237 17918 8265
rect 18201 8237 18302 8265
rect 20674 8191 20702 8339
rect 21442 8311 21950 8339
rect 22978 8311 23294 8339
rect 23362 8311 23390 8385
rect 23481 8311 23568 8339
rect 25474 8311 25598 8339
rect 23746 8237 25310 8265
rect 23746 8191 23774 8237
rect 18082 8163 20702 8191
rect 21730 8163 23774 8191
rect 25282 8191 25310 8237
rect 25282 8163 28574 8191
rect 3298 8089 3518 8117
rect 8578 8089 8702 8117
rect 9154 8089 9278 8117
rect 14722 8089 16670 8117
rect 22114 8089 22238 8117
rect 24226 8089 24350 8117
rect 25378 8089 25502 8117
rect 0 7943 32064 8041
rect 1666 7867 1886 7895
rect 2626 7867 3134 7895
rect 7234 7867 7358 7895
rect 10905 7867 10992 7895
rect 11746 7867 13022 7895
rect 14146 7867 14366 7895
rect 9922 7793 11678 7821
rect 11746 7747 11774 7867
rect 14338 7821 14366 7867
rect 14818 7867 15038 7895
rect 15394 7867 16478 7895
rect 14818 7821 14846 7867
rect 11938 7793 12542 7821
rect 14338 7793 14846 7821
rect 15202 7793 15326 7821
rect 12514 7784 12542 7793
rect 12514 7756 13118 7784
rect 706 7719 1406 7747
rect 1858 7719 2942 7747
rect 3106 7719 3326 7747
rect 4738 7719 4958 7747
rect 7042 7719 7166 7747
rect 7234 7719 7358 7747
rect 8674 7719 9854 7747
rect 10882 7719 11006 7747
rect 11673 7719 11774 7747
rect 13090 7747 13118 7756
rect 13090 7719 13694 7747
rect 7234 7673 7262 7719
rect 10882 7673 10910 7719
rect 4258 7645 4478 7673
rect 4546 7645 5534 7673
rect 6850 7645 7262 7673
rect 9922 7645 10910 7673
rect 11842 7645 11966 7673
rect 12322 7645 12830 7673
rect 12921 7645 13008 7673
rect 13762 7645 14078 7673
rect 14146 7645 14750 7673
rect 15298 7645 15326 7793
rect 16450 7719 16478 7867
rect 21058 7793 21566 7821
rect 16569 7719 16656 7747
rect 20098 7719 20318 7747
rect 20482 7719 20702 7747
rect 21442 7719 22142 7747
rect 21561 7645 21648 7673
rect 21730 7645 21854 7673
rect 21922 7645 22814 7673
rect 14242 7571 15518 7599
rect 16834 7571 17438 7599
rect 16834 7525 16862 7571
rect 1666 7497 2942 7525
rect 1666 7451 1694 7497
rect 1474 7423 1694 7451
rect 2914 7451 2942 7497
rect 16450 7497 16862 7525
rect 16450 7451 16478 7497
rect 2914 7423 3134 7451
rect 4066 7423 4478 7451
rect 10329 7423 10416 7451
rect 11938 7423 12158 7451
rect 12994 7423 13310 7451
rect 13762 7423 14078 7451
rect 14530 7423 15134 7451
rect 15202 7423 16478 7451
rect 17410 7451 17438 7571
rect 19330 7571 19934 7599
rect 19330 7451 19358 7571
rect 19906 7525 19934 7571
rect 19906 7497 20222 7525
rect 17410 7423 17630 7451
rect 19138 7423 19358 7451
rect 20194 7451 20222 7497
rect 20194 7423 20414 7451
rect 0 7277 32064 7375
rect 610 7201 734 7229
rect 1017 7201 1104 7229
rect 2146 7201 2654 7229
rect 2626 7081 2654 7201
rect 3490 7201 3998 7229
rect 5122 7201 5438 7229
rect 5506 7201 6110 7229
rect 9154 7201 9470 7229
rect 10329 7201 10416 7229
rect 11458 7201 11774 7229
rect 13186 7201 13790 7229
rect 14265 7201 14352 7229
rect 14434 7201 15230 7229
rect 17721 7201 17808 7229
rect 22786 7201 23006 7229
rect 26722 7201 26942 7229
rect 3490 7081 3518 7201
rect 26914 7155 26942 7201
rect 27394 7201 27614 7229
rect 27394 7155 27422 7201
rect 7042 7127 8510 7155
rect 26914 7127 27422 7155
rect 1474 7053 1886 7081
rect 2338 7053 2462 7081
rect 2626 7053 3518 7081
rect 3874 7053 4094 7081
rect 10594 7053 11102 7081
rect 1474 7007 1502 7053
rect 802 6979 1502 7007
rect 1689 6979 1776 7007
rect 1858 6979 1886 7053
rect 10594 7007 10622 7053
rect 3682 6979 3902 7007
rect 4930 6979 5342 7007
rect 5890 6979 6014 7007
rect 7234 6979 7358 7007
rect 7330 6933 7358 6979
rect 8194 6979 9086 7007
rect 9177 6979 9264 7007
rect 9730 6979 10334 7007
rect 10402 6979 10622 7007
rect 11074 7007 11102 7053
rect 15778 7053 17150 7081
rect 19042 7053 19166 7081
rect 25401 7053 25488 7081
rect 15778 7007 15806 7053
rect 11074 6979 11294 7007
rect 11554 6979 11870 7007
rect 13017 6979 13104 7007
rect 610 6905 734 6933
rect 898 6859 926 6933
rect 1570 6905 2270 6933
rect 7330 6905 8126 6933
rect 1570 6859 1598 6905
rect 8194 6859 8222 6979
rect 10402 6933 10430 6979
rect 10018 6905 10430 6933
rect 12322 6905 12926 6933
rect 13186 6859 13214 7007
rect 13282 6979 14270 7007
rect 15394 6979 15806 7007
rect 17122 7007 17150 7053
rect 17122 6979 17342 7007
rect 17698 6979 19550 7007
rect 23170 6979 24350 7007
rect 24418 6979 25406 7007
rect 27120 6979 27710 7007
rect 13977 6905 14064 6933
rect 15874 6905 16190 6933
rect 16354 6905 17630 6933
rect 22905 6905 22992 6933
rect 23074 6905 23294 6933
rect 25186 6905 25790 6933
rect 226 6831 1598 6859
rect 8098 6831 8222 6859
rect 10594 6831 12158 6859
rect 8098 6785 8126 6831
rect 12130 6822 12158 6831
rect 12802 6831 13214 6859
rect 12802 6822 12830 6831
rect 12130 6794 12830 6822
rect 2073 6757 2160 6785
rect 5026 6757 5630 6785
rect 7234 6757 8126 6785
rect 8194 6757 8318 6785
rect 16281 6757 16368 6785
rect 19330 6757 19742 6785
rect 24130 6757 24446 6785
rect 0 6611 32064 6709
rect 2338 6535 3038 6563
rect 3490 6535 4286 6563
rect 4354 6535 4958 6563
rect 7138 6535 7262 6563
rect 13378 6535 13790 6563
rect 13762 6526 13790 6535
rect 14338 6535 14558 6563
rect 15394 6535 15614 6563
rect 17602 6535 17726 6563
rect 21826 6535 21950 6563
rect 22306 6535 23102 6563
rect 25378 6535 25502 6563
rect 14338 6526 14366 6535
rect 13762 6498 14366 6526
rect 4546 6461 6014 6489
rect 7906 6461 8510 6489
rect 7906 6415 7934 6461
rect 1954 6387 2270 6415
rect 2242 6341 2270 6387
rect 3010 6387 3230 6415
rect 3298 6387 4766 6415
rect 5817 6387 5904 6415
rect 6105 6387 6192 6415
rect 7714 6387 7934 6415
rect 8482 6415 8510 6461
rect 10786 6461 13598 6489
rect 10786 6415 10814 6461
rect 8482 6387 8702 6415
rect 8770 6387 10814 6415
rect 13570 6415 13598 6461
rect 13570 6387 14558 6415
rect 19714 6387 19838 6415
rect 20578 6387 20702 6415
rect 23074 6387 23198 6415
rect 3010 6341 3038 6387
rect 2242 6313 3038 6341
rect 3202 6313 3230 6387
rect 8770 6341 8798 6387
rect 4450 6313 4574 6341
rect 4930 6313 5150 6341
rect 4450 6267 4478 6313
rect 3394 6239 4478 6267
rect 5122 6267 5150 6313
rect 5890 6313 6110 6341
rect 6370 6313 6878 6341
rect 8025 6313 8798 6341
rect 9250 6313 9470 6341
rect 5890 6267 5918 6313
rect 5122 6239 5918 6267
rect 9250 6253 9278 6313
rect 9442 6267 9470 6313
rect 10114 6313 10512 6341
rect 11952 6313 12638 6341
rect 10114 6267 10142 6313
rect 12610 6267 12638 6313
rect 13474 6313 13680 6341
rect 15120 6313 15902 6341
rect 19353 6313 19440 6341
rect 20098 6313 20510 6341
rect 20578 6313 20606 6387
rect 23266 6341 23294 6415
rect 23650 6387 26270 6415
rect 20674 6313 20798 6341
rect 21058 6313 23294 6341
rect 24345 6313 24432 6341
rect 26434 6313 26942 6341
rect 13474 6267 13502 6313
rect 9442 6239 10142 6267
rect 10306 6239 11102 6267
rect 12610 6239 13502 6267
rect 15874 6267 15902 6313
rect 15874 6239 18288 6267
rect 20674 6193 20702 6313
rect 29314 6239 31742 6267
rect 11746 6165 12254 6193
rect 19138 6165 20702 6193
rect 21154 6165 22142 6193
rect 11746 6119 11774 6165
rect 9250 6091 9950 6119
rect 11554 6091 11774 6119
rect 12226 6119 12254 6165
rect 21154 6119 21182 6165
rect 12226 6091 12446 6119
rect 20962 6091 21182 6119
rect 22114 6119 22142 6165
rect 29314 6119 29342 6239
rect 22114 6091 22334 6119
rect 23458 6091 24542 6119
rect 26626 6091 26846 6119
rect 29122 6091 29342 6119
rect 31714 6119 31742 6239
rect 31714 6091 31934 6119
rect 0 5945 32064 6043
rect 610 5869 734 5897
rect 4834 5869 4958 5897
rect 6178 5869 6398 5897
rect 11842 5869 11966 5897
rect 13017 5869 13104 5897
rect 14722 5869 15326 5897
rect 15874 5869 16670 5897
rect 20025 5869 20112 5897
rect 24322 5869 24926 5897
rect 28738 5869 28958 5897
rect 5794 5795 6686 5823
rect 22114 5795 22910 5823
rect 1282 5721 1790 5749
rect 4066 5721 4286 5749
rect 8194 5721 8318 5749
rect 12130 5721 12734 5749
rect 1282 5675 1310 5721
rect 130 5647 1310 5675
rect 1762 5675 1790 5721
rect 4162 5675 4190 5721
rect 12130 5675 12158 5721
rect 1762 5647 1982 5675
rect 3874 5647 3998 5675
rect 1954 5601 1982 5647
rect 4066 5601 4094 5675
rect 4162 5647 4574 5675
rect 5721 5647 5808 5675
rect 9177 5647 9264 5675
rect 10306 5647 10430 5675
rect 10498 5647 10622 5675
rect 11481 5647 11568 5675
rect 1401 5573 1488 5601
rect 1954 5573 2366 5601
rect 2722 5573 2942 5601
rect 3033 5573 3120 5601
rect 3202 5573 4094 5601
rect 8002 5573 8222 5601
rect 11650 5527 11678 5675
rect 11746 5647 12158 5675
rect 12706 5675 12734 5721
rect 19618 5721 20784 5749
rect 22114 5735 22142 5795
rect 22233 5721 22320 5749
rect 22882 5735 22910 5795
rect 24226 5795 24446 5823
rect 24226 5735 24254 5795
rect 24418 5786 24446 5795
rect 24994 5795 26942 5823
rect 24994 5786 25022 5795
rect 24418 5758 25022 5786
rect 26914 5749 26942 5795
rect 27490 5795 27710 5823
rect 27490 5749 27518 5795
rect 12706 5647 13022 5675
rect 13858 5647 14078 5675
rect 16354 5647 16478 5675
rect 16752 5647 16839 5675
rect 17314 5647 18192 5675
rect 19618 5661 19646 5721
rect 25378 5675 25406 5749
rect 26914 5721 27518 5749
rect 28930 5749 28958 5869
rect 31810 5869 32030 5897
rect 31810 5749 31838 5869
rect 28930 5721 31838 5749
rect 21730 5647 23294 5675
rect 21730 5601 21758 5647
rect 23266 5601 23294 5647
rect 24994 5647 25214 5675
rect 25378 5647 25598 5675
rect 24994 5601 25022 5647
rect 15394 5573 15806 5601
rect 19426 5573 19646 5601
rect 19714 5573 19838 5601
rect 19906 5573 21758 5601
rect 22690 5573 22814 5601
rect 23266 5573 25022 5601
rect 25570 5601 25598 5647
rect 26146 5647 26558 5675
rect 26146 5601 26174 5647
rect 25570 5573 26174 5601
rect 26361 5573 26448 5601
rect 26626 5573 26750 5601
rect 19618 5527 19646 5573
rect 19906 5527 19934 5573
rect 10882 5499 11678 5527
rect 12034 5499 13310 5527
rect 19618 5499 19934 5527
rect 1474 5425 1598 5453
rect 3106 5425 3902 5453
rect 8578 5425 8990 5453
rect 10402 5425 10718 5453
rect 14146 5425 14270 5453
rect 15033 5425 15120 5453
rect 16185 5425 16272 5453
rect 17625 5425 17712 5453
rect 26626 5425 26750 5453
rect 0 5279 32064 5377
rect 2146 5203 3230 5231
rect 3874 5203 4190 5231
rect 8578 5203 8702 5231
rect 11001 5203 11088 5231
rect 12825 5203 12912 5231
rect 13666 5203 14078 5231
rect 16738 5203 17438 5231
rect 19618 5203 19742 5231
rect 20985 5203 21072 5231
rect 22786 5203 23006 5231
rect 24153 5203 24240 5231
rect 26242 5203 26462 5231
rect 26434 5157 26462 5203
rect 27586 5203 28094 5231
rect 27586 5157 27614 5203
rect 2626 5129 3038 5157
rect 3394 5129 3614 5157
rect 5794 5129 6014 5157
rect 7138 5129 10814 5157
rect 23074 5129 24446 5157
rect 26434 5129 27614 5157
rect 28066 5157 28094 5203
rect 29506 5203 29726 5231
rect 29506 5157 29534 5203
rect 28066 5129 29534 5157
rect 2338 4981 2942 5009
rect 3010 4981 3038 5129
rect 3225 5055 3312 5083
rect 3586 5009 3614 5129
rect 4258 5055 4574 5083
rect 4834 5055 5534 5083
rect 4258 5009 4286 5055
rect 3586 4981 4286 5009
rect 5122 4981 5246 5009
rect 5506 4981 5534 5055
rect 5794 5055 6686 5083
rect 5794 4981 5822 5055
rect 5890 4981 6014 5009
rect 7138 4981 7166 5129
rect 23074 5083 23102 5129
rect 8674 5055 8798 5083
rect 10690 5055 11198 5083
rect 12802 5055 13406 5083
rect 13474 5055 13598 5083
rect 15202 5055 16286 5083
rect 18178 5055 19070 5083
rect 13474 5009 13502 5055
rect 18178 5009 18206 5055
rect 7522 4981 8318 5009
rect 8482 4981 8606 5009
rect 10594 4981 11006 5009
rect 12130 4981 12350 5009
rect 12898 4981 13502 5009
rect 14530 4981 15614 5009
rect 17698 4981 18206 5009
rect 19042 5009 19070 5055
rect 19234 5009 19262 5083
rect 22882 5055 23102 5083
rect 27801 5055 27888 5083
rect 19042 4981 19358 5009
rect 20098 4981 21086 5009
rect 21168 4981 21255 5009
rect 21346 4981 21470 5009
rect 23074 4981 24254 5009
rect 4450 4907 5054 4935
rect 5026 4861 5054 4907
rect 5890 4861 5918 4981
rect 7522 4935 7550 4981
rect 7042 4907 7550 4935
rect 8290 4935 8318 4981
rect 24226 4935 24254 4981
rect 24418 4981 24542 5009
rect 26722 4981 26942 5009
rect 24418 4935 24446 4981
rect 8290 4907 9566 4935
rect 16752 4907 17342 4935
rect 19234 4907 19358 4935
rect 24226 4907 24446 4935
rect 26914 4935 26942 4981
rect 27394 4981 27614 5009
rect 27682 4981 27792 5009
rect 27394 4935 27422 4981
rect 26914 4907 27422 4935
rect 5026 4833 5918 4861
rect 7618 4833 9950 4861
rect 11170 4833 11678 4861
rect 11170 4787 11198 4833
rect 6873 4759 6960 4787
rect 8290 4759 9182 4787
rect 10882 4759 11198 4787
rect 11650 4787 11678 4833
rect 18274 4833 19070 4861
rect 18274 4787 18302 4833
rect 11650 4759 11870 4787
rect 18082 4759 18302 4787
rect 19042 4787 19070 4833
rect 19522 4833 20606 4861
rect 19522 4787 19550 4833
rect 19042 4759 19550 4787
rect 20578 4787 20606 4833
rect 20578 4759 20798 4787
rect 0 4613 32064 4711
rect 1474 4537 1886 4565
rect 2722 4537 2846 4565
rect 8770 4537 9182 4565
rect 12249 4537 12336 4565
rect 16738 4537 16958 4565
rect 10978 4500 11678 4528
rect 10978 4491 11006 4500
rect 10786 4463 11006 4491
rect 11650 4491 11678 4500
rect 16930 4491 16958 4537
rect 17794 4537 18302 4565
rect 20386 4537 20702 4565
rect 21442 4537 21758 4565
rect 23458 4537 23678 4565
rect 11650 4463 11870 4491
rect 8386 4426 9182 4454
rect 8386 4417 8414 4426
rect 2242 4389 2846 4417
rect 2914 4389 3134 4417
rect 8194 4389 8414 4417
rect 9154 4417 9182 4426
rect 9154 4389 9374 4417
rect 9346 4343 9374 4389
rect 11842 4343 11870 4463
rect 12706 4463 13214 4491
rect 16930 4463 17150 4491
rect 12706 4343 12734 4463
rect 17122 4417 17150 4463
rect 17794 4417 17822 4537
rect 23650 4491 23678 4537
rect 24130 4537 24350 4565
rect 26242 4537 26462 4565
rect 24130 4491 24158 4537
rect 18009 4463 18096 4491
rect 23650 4463 24158 4491
rect 17122 4389 17822 4417
rect 130 4315 542 4343
rect 1474 4315 2078 4343
rect 2146 4269 2174 4343
rect 2914 4315 3038 4343
rect 3490 4315 3710 4343
rect 8578 4315 9086 4343
rect 9154 4315 9278 4343
rect 9346 4315 10526 4343
rect 11842 4315 12734 4343
rect 12898 4315 13406 4343
rect 14434 4315 15422 4343
rect 15778 4315 16766 4343
rect 18178 4315 19166 4343
rect 13378 4269 13406 4315
rect 16738 4269 16766 4315
rect 19138 4269 19166 4315
rect 20674 4315 21662 4343
rect 20674 4269 20702 4315
rect 26242 4269 26270 4537
rect 26434 4528 26462 4537
rect 28546 4537 28766 4565
rect 28546 4528 28574 4537
rect 26434 4500 28574 4528
rect 26530 4389 28670 4417
rect 28738 4343 28766 4537
rect 28450 4269 28478 4343
rect 28738 4315 29630 4343
rect 994 4241 1406 4269
rect 1378 4195 1406 4241
rect 1954 4241 2462 4269
rect 10114 4241 11006 4269
rect 13378 4241 13502 4269
rect 14242 4241 14654 4269
rect 16450 4241 16670 4269
rect 16738 4241 16862 4269
rect 18850 4241 19070 4269
rect 19138 4241 19262 4269
rect 19810 4241 20702 4269
rect 23650 4241 24254 4269
rect 24418 4241 24542 4269
rect 26146 4241 26270 4269
rect 27202 4241 28478 4269
rect 1954 4195 1982 4241
rect 27202 4195 27230 4241
rect 1378 4167 1982 4195
rect 3970 4167 4478 4195
rect 3970 4121 3998 4167
rect 3778 4093 3998 4121
rect 4450 4121 4478 4167
rect 26434 4167 27230 4195
rect 26434 4121 26462 4167
rect 4450 4093 4670 4121
rect 13474 4093 14270 4121
rect 14530 4093 14846 4121
rect 18274 4093 19262 4121
rect 20866 4093 21086 4121
rect 25954 4093 26462 4121
rect 28185 4093 28272 4121
rect 0 3947 32064 4045
rect 3010 3871 3134 3899
rect 4738 3871 5150 3899
rect 9657 3871 9744 3899
rect 16761 3871 16848 3899
rect 18562 3871 18686 3899
rect 19737 3871 19824 3899
rect 24514 3871 24734 3899
rect 24706 3825 24734 3871
rect 25570 3871 25790 3899
rect 25570 3825 25598 3871
rect 14626 3797 16574 3825
rect 14914 3751 14942 3797
rect 16546 3751 16574 3797
rect 17890 3797 18302 3825
rect 17890 3751 17918 3797
rect 18274 3788 18302 3797
rect 18754 3797 19454 3825
rect 20578 3797 21278 3825
rect 21442 3797 22910 3825
rect 24706 3797 25598 3825
rect 26073 3797 26160 3825
rect 18754 3788 18782 3797
rect 18274 3760 18782 3788
rect 20578 3751 20606 3797
rect 1570 3723 2750 3751
rect 2818 3723 3038 3751
rect 4642 3723 5246 3751
rect 6946 3723 7646 3751
rect 7833 3723 7920 3751
rect 14722 3723 14846 3751
rect 14914 3723 15038 3751
rect 16546 3723 17918 3751
rect 20386 3723 20606 3751
rect 21250 3751 21278 3797
rect 21250 3723 21662 3751
rect 2434 3649 2942 3677
rect 3010 3649 3038 3723
rect 5218 3677 5246 3723
rect 5218 3649 5918 3677
rect 6082 3649 6206 3677
rect 9264 3649 14928 3677
rect 18178 3649 18302 3677
rect 18370 3649 19358 3677
rect 19426 3649 20304 3677
rect 22114 3649 22622 3677
rect 23097 3649 24638 3677
rect 322 3575 1406 3603
rect 322 3529 350 3575
rect 130 3501 350 3529
rect 1378 3529 1406 3575
rect 3202 3575 4286 3603
rect 3202 3529 3230 3575
rect 1378 3501 3230 3529
rect 4258 3529 4286 3575
rect 19330 3529 19358 3649
rect 22114 3603 22142 3649
rect 21922 3575 22142 3603
rect 22594 3603 22622 3649
rect 24610 3603 24638 3649
rect 25666 3649 25982 3677
rect 25666 3603 25694 3649
rect 22594 3575 22814 3603
rect 24610 3575 25694 3603
rect 4258 3501 4574 3529
rect 19330 3501 21758 3529
rect 21730 3492 21758 3501
rect 21730 3464 22526 3492
rect 22498 3455 22526 3464
rect 6082 3427 6878 3455
rect 17890 3427 18014 3455
rect 22498 3427 23102 3455
rect 0 3281 32064 3379
rect 3298 3205 3518 3233
rect 3490 3159 3518 3205
rect 4066 3205 4286 3233
rect 6585 3205 6672 3233
rect 10978 3205 11102 3233
rect 13017 3205 13104 3233
rect 16450 3205 16574 3233
rect 18658 3205 18878 3233
rect 4066 3159 4094 3205
rect 18850 3159 18878 3205
rect 19714 3205 19934 3233
rect 20962 3205 21182 3233
rect 22713 3205 22800 3233
rect 19714 3159 19742 3205
rect 22978 3159 23006 3233
rect 23097 3205 23184 3233
rect 24610 3205 24734 3233
rect 29529 3205 29616 3233
rect 3490 3131 4094 3159
rect 4354 3131 5342 3159
rect 18850 3131 19742 3159
rect 22617 3131 22704 3159
rect 22978 3131 24446 3159
rect 4354 3011 4382 3131
rect 17794 3057 17918 3085
rect 27490 3057 28286 3085
rect 3106 2983 4382 3011
rect 4450 2983 6110 3011
rect 10809 2983 10896 3011
rect 12706 2983 13022 3011
rect 13282 2983 13886 3011
rect 15778 2983 16478 3011
rect 21081 2983 21168 3011
rect 21442 2983 23006 3011
rect 23650 2983 24350 3011
rect 27010 2983 27696 3011
rect 5506 2909 5630 2937
rect 6585 2909 6672 2937
rect 6777 2909 6864 2937
rect 8770 2909 8990 2937
rect 9058 2909 9950 2937
rect 10690 2909 11102 2937
rect 18009 2909 18302 2937
rect 5506 2863 5534 2909
rect 18274 2863 18302 2909
rect 19522 2909 20414 2937
rect 26818 2909 27038 2937
rect 19522 2863 19550 2909
rect 3490 2835 5534 2863
rect 5602 2835 6782 2863
rect 14050 2835 14558 2863
rect 18274 2835 19550 2863
rect 27010 2863 27038 2909
rect 27586 2909 27902 2937
rect 30274 2909 31934 2937
rect 27586 2863 27614 2909
rect 27010 2835 27614 2863
rect 9346 2798 10526 2826
rect 9346 2789 9374 2798
rect 9081 2761 9374 2789
rect 10498 2789 10526 2798
rect 14050 2789 14078 2835
rect 10498 2761 10718 2789
rect 13474 2761 14078 2789
rect 14530 2789 14558 2835
rect 14530 2761 14750 2789
rect 0 2615 32064 2713
rect 5602 2539 5918 2567
rect 6082 2539 6302 2567
rect 10617 2539 10704 2567
rect 10809 2539 10896 2567
rect 12633 2539 12720 2567
rect 15202 2539 15806 2567
rect 21154 2539 21374 2567
rect 5602 2493 5630 2539
rect 21346 2530 21374 2539
rect 22018 2539 22238 2567
rect 27106 2539 27422 2567
rect 22018 2530 22046 2539
rect 21346 2502 22046 2530
rect 3394 2465 5630 2493
rect 14626 2465 15518 2493
rect 2914 2391 3134 2419
rect 3394 2345 3422 2465
rect 14626 2419 14654 2465
rect 4546 2391 4766 2419
rect 4738 2345 4766 2391
rect 5698 2391 5918 2419
rect 8674 2391 10526 2419
rect 14457 2391 14654 2419
rect 14722 2391 14846 2419
rect 3298 2317 3422 2345
rect 4066 2317 4478 2345
rect 4738 2317 5150 2345
rect 4066 2271 4094 2317
rect 2722 2243 4094 2271
rect 5122 2271 5150 2317
rect 5698 2271 5726 2391
rect 8674 2345 8702 2391
rect 15490 2345 15518 2465
rect 27394 2419 27422 2539
rect 31810 2539 32030 2567
rect 31810 2419 31838 2539
rect 15970 2391 16862 2419
rect 15970 2345 15998 2391
rect 5986 2317 6110 2345
rect 6192 2317 6279 2345
rect 8578 2317 8702 2345
rect 8793 2317 8880 2345
rect 14626 2271 14654 2331
rect 15490 2317 15998 2345
rect 16834 2345 16862 2391
rect 17314 2391 18302 2419
rect 16834 2317 17054 2345
rect 17314 2271 17342 2391
rect 18274 2345 18302 2391
rect 21154 2391 21662 2419
rect 21154 2345 21182 2391
rect 18274 2317 20222 2345
rect 20313 2317 21182 2345
rect 21634 2345 21662 2391
rect 23842 2391 24926 2419
rect 23842 2345 23870 2391
rect 21634 2317 23870 2345
rect 24898 2345 24926 2391
rect 25570 2391 26558 2419
rect 27394 2391 31838 2419
rect 25570 2345 25598 2391
rect 24898 2317 25598 2345
rect 26530 2345 26558 2391
rect 26530 2317 26846 2345
rect 5122 2243 5726 2271
rect 7234 2243 8222 2271
rect 8674 2243 8798 2271
rect 14626 2243 15888 2271
rect 17232 2243 17342 2271
rect 17410 2243 18206 2271
rect 20002 2243 20126 2271
rect 20194 2257 20222 2317
rect 27106 2243 27230 2271
rect 3298 2169 3518 2197
rect 7234 2123 7262 2243
rect 4857 2095 4944 2123
rect 7042 2095 7262 2123
rect 8194 2123 8222 2243
rect 23938 2169 24830 2197
rect 23938 2123 23966 2169
rect 8194 2095 8414 2123
rect 23746 2095 23966 2123
rect 24802 2123 24830 2169
rect 24802 2095 25022 2123
rect 0 1949 32064 2047
rect 3106 1873 3230 1901
rect 6082 1873 6206 1901
rect 6658 1827 6686 1901
rect 8866 1873 9182 1901
rect 20098 1873 20894 1901
rect 24322 1873 24542 1901
rect 5794 1799 6686 1827
rect 10306 1753 10334 1827
rect 20674 1799 20798 1827
rect 24514 1753 24542 1873
rect 26914 1873 27134 1901
rect 26914 1753 26942 1873
rect 4546 1725 5726 1753
rect 6946 1725 7070 1753
rect 8496 1725 10416 1753
rect 12322 1725 13022 1753
rect 13186 1725 14462 1753
rect 23458 1725 23966 1753
rect 24514 1725 26942 1753
rect 5698 1679 5726 1725
rect 34 1651 2846 1679
rect 3321 1651 3408 1679
rect 5602 1605 5630 1679
rect 5698 1651 6110 1679
rect 6178 1651 6302 1679
rect 7330 1651 8126 1679
rect 6178 1605 6206 1651
rect 5602 1577 6206 1605
rect 8098 1605 8126 1651
rect 10018 1651 10622 1679
rect 10018 1605 10046 1651
rect 12322 1605 12350 1725
rect 8098 1577 10046 1605
rect 10210 1577 12350 1605
rect 12994 1605 13022 1725
rect 14553 1651 14640 1679
rect 20985 1651 21072 1679
rect 23650 1651 23870 1679
rect 24057 1651 24144 1679
rect 12994 1577 14846 1605
rect 21154 1577 21278 1605
rect 12610 1466 13310 1494
rect 12610 1457 12638 1466
rect 12418 1429 12638 1457
rect 13282 1457 13310 1466
rect 13282 1429 14270 1457
rect 0 1283 32064 1381
rect 4761 1207 4848 1235
rect 13401 1207 13488 1235
rect 15586 1207 16670 1235
rect 18105 1207 18192 1235
rect 20674 1207 20990 1235
rect 16642 1161 16670 1207
rect 10690 1059 13214 1087
rect 16450 1013 16478 1161
rect 16642 1133 17918 1161
rect 17890 1087 17918 1133
rect 17890 1059 18302 1087
rect 23385 1059 23472 1087
rect 23577 1059 23664 1087
rect 130 985 3326 1013
rect 3682 985 4478 1013
rect 4546 985 4958 1013
rect 13282 985 15902 1013
rect 15970 985 18110 1013
rect 20866 985 20990 1013
rect 21058 985 24158 1013
rect 3298 911 3614 939
rect 15874 865 15902 985
rect 15874 837 17918 865
rect 0 617 32064 715
rect 0 -49 32064 49
<< metal2 >>
rect 31967 32583 32064 32611
rect 0 32509 97 32537
rect 34 32361 62 32509
rect 0 31177 97 31205
rect 2050 31177 2078 31649
rect 34 31103 62 31177
rect 3106 30909 3134 31057
rect 3010 30881 3134 30909
rect 3010 30391 3038 30881
rect 3010 30363 3134 30391
rect 0 29845 97 29873
rect 2050 29845 2078 30243
rect 34 29475 62 29845
rect 1954 29133 1982 29577
rect 1858 29105 1982 29133
rect 0 28439 158 28467
rect 1858 28245 1886 29105
rect 2146 28291 2174 29651
rect 1858 28217 1982 28245
rect 1954 28097 1982 28217
rect 1954 28069 2174 28097
rect 34 27135 62 27727
rect 1282 27551 1502 27579
rect 0 27107 97 27135
rect 34 25803 62 26469
rect 0 25775 97 25803
rect 34 24397 62 25581
rect 802 24517 830 25655
rect 0 24369 97 24397
rect 1282 23629 1310 27551
rect 1954 27181 1982 28069
rect 1666 24101 1694 24767
rect 1474 24073 1694 24101
rect 1474 23851 1502 24073
rect 0 23037 97 23065
rect 34 22889 62 23037
rect 34 21733 62 21807
rect 0 21705 97 21733
rect 1186 20521 1214 21585
rect 0 20373 97 20401
rect 34 20151 62 20373
rect 226 20105 254 20475
rect 1378 20299 1406 20771
rect 1570 20521 1598 21067
rect 34 20077 254 20105
rect 34 18995 62 20077
rect 0 18967 97 18995
rect 994 17857 1022 18329
rect 2050 17709 2078 21733
rect 2434 21705 2462 27061
rect 0 17635 97 17663
rect 34 16377 62 17635
rect 0 16303 97 16331
rect 34 16155 62 16303
rect 34 14925 62 15073
rect 0 14897 97 14925
rect 34 13593 62 14259
rect 0 13565 97 13593
rect 226 13519 254 16775
rect 2722 16525 2750 29651
rect 3106 29577 3134 30363
rect 3298 29651 3326 30983
rect 4162 30909 4190 31649
rect 4162 30881 4286 30909
rect 3298 29623 3422 29651
rect 3010 29549 3134 29577
rect 3010 28837 3038 29549
rect 3010 28809 3134 28837
rect 3106 28467 3134 28809
rect 3010 28439 3134 28467
rect 3010 27505 3038 28439
rect 3010 27477 3134 27505
rect 3106 27033 3134 27477
rect 3298 25507 3326 29577
rect 4258 27625 4286 30881
rect 4738 27625 4766 30095
rect 5506 27579 5534 29799
rect 5986 28513 6014 29651
rect 6274 28911 6302 31427
rect 6562 30955 6590 31575
rect 6754 28957 6782 31427
rect 8290 30909 8318 31427
rect 8290 30881 8414 30909
rect 7426 29697 7454 30761
rect 8098 29577 8126 29725
rect 6274 28883 6686 28911
rect 6178 27653 6206 28319
rect 6658 27847 6686 28883
rect 6082 27625 6206 27653
rect 3490 26737 3518 27431
rect 3874 26293 3902 26765
rect 3298 25479 3422 25507
rect 3106 24961 3134 25433
rect 3394 24915 3422 25479
rect 4258 25063 4286 27431
rect 3298 24887 3422 24915
rect 4162 25035 4286 25063
rect 2914 23435 2942 24101
rect 2914 23407 3134 23435
rect 2914 22519 2942 23139
rect 3106 21187 3134 23407
rect 3298 23065 3326 24887
rect 4162 24175 4190 25035
rect 4450 24221 4478 27579
rect 5506 27551 5726 27579
rect 4642 27357 4670 27505
rect 4642 27329 4766 27357
rect 4738 26765 4766 27329
rect 4642 26737 4766 26765
rect 4642 25035 4670 26737
rect 5026 26617 5054 26765
rect 4930 26589 5054 26617
rect 4930 25109 4958 26589
rect 5506 26219 5534 27551
rect 6082 27135 6110 27625
rect 6370 27181 6398 27579
rect 6082 27107 6206 27135
rect 6178 25849 6206 27107
rect 7522 26959 7550 29577
rect 8002 29549 8126 29577
rect 8002 28985 8030 29549
rect 8002 28957 8126 28985
rect 8290 28957 8318 30881
rect 8674 30511 8702 31649
rect 9538 30881 9566 31649
rect 7906 28467 7934 28763
rect 7810 28439 7934 28467
rect 7810 27801 7838 28439
rect 7810 27773 7934 27801
rect 7906 27625 7934 27773
rect 8098 27357 8126 28957
rect 8482 27875 8510 30095
rect 9730 29059 9758 30317
rect 11842 29651 11870 29799
rect 11650 29623 11870 29651
rect 12322 29623 12350 31649
rect 9538 29031 9758 29059
rect 9538 28467 9566 29031
rect 9538 28439 9662 28467
rect 8482 27847 8702 27875
rect 8482 27727 8510 27847
rect 9250 27801 9278 28097
rect 9154 27773 9278 27801
rect 8482 27699 8606 27727
rect 8002 27329 8126 27357
rect 8002 27209 8030 27329
rect 7810 27181 8030 27209
rect 4162 24147 4286 24175
rect 3250 23037 3326 23065
rect 3250 22473 3278 23037
rect 3394 22519 3422 22991
rect 3250 22445 3326 22473
rect 3298 21779 3326 22445
rect 3106 19559 3134 20771
rect 3298 20299 3326 21437
rect 3874 21215 3902 23657
rect 4258 22473 4286 24147
rect 4354 23703 4382 24101
rect 4162 22445 4286 22473
rect 4162 21511 4190 22445
rect 4450 21557 4478 22991
rect 4546 22963 4574 24175
rect 5602 23879 5630 24249
rect 5602 23851 5726 23879
rect 5602 23805 5630 23851
rect 5506 23777 5630 23805
rect 4738 22177 4766 23435
rect 5506 23213 5534 23777
rect 5794 23703 5822 24767
rect 5986 24517 6014 25063
rect 5410 23185 5534 23213
rect 5410 22371 5438 23185
rect 5794 23065 5822 23583
rect 5698 23037 5822 23065
rect 5986 23407 6110 23435
rect 5698 22547 5726 23037
rect 5698 22519 5822 22547
rect 5794 22371 5822 22519
rect 4738 22149 4862 22177
rect 4162 21483 4286 21511
rect 3874 21187 3998 21215
rect 3970 20151 3998 21187
rect 4162 20447 4190 20771
rect 4258 19735 4286 21483
rect 3298 19041 3326 19439
rect 3682 19291 3710 19439
rect 3586 19263 3710 19291
rect 3586 18255 3614 19263
rect 3874 18773 3902 19735
rect 4162 19707 4286 19735
rect 4162 18921 4190 19707
rect 4162 18893 4286 18921
rect 3778 18745 3902 18773
rect 3874 18301 3902 18745
rect 4258 18551 4286 18893
rect 4162 18523 4286 18551
rect 4162 18375 4190 18523
rect 4354 18449 4382 19661
rect 3586 18227 3710 18255
rect 3298 17663 3326 18107
rect 3298 17635 3422 17663
rect 3682 17635 3710 18227
rect 3202 17191 3230 17589
rect 3394 17145 3422 17635
rect 3298 17117 3422 17145
rect 3298 16969 3326 17117
rect 706 13639 734 15147
rect 1186 13593 1214 13741
rect 34 13491 254 13519
rect 994 13565 1214 13593
rect 34 12261 62 13491
rect 0 12233 97 12261
rect 34 10855 62 11003
rect 0 10827 97 10855
rect 130 10781 158 12409
rect 610 11567 638 12335
rect 994 12261 1022 13565
rect 1378 13445 1406 14925
rect 2146 13861 2174 14999
rect 2434 13741 2462 16331
rect 3106 15193 3134 15665
rect 3394 15147 3422 16109
rect 3394 15119 3518 15147
rect 2626 14703 2654 14851
rect 2626 14675 2750 14703
rect 2722 14185 2750 14675
rect 2338 13713 2462 13741
rect 2626 14157 2750 14185
rect 1282 13417 1406 13445
rect 1282 12483 1310 13417
rect 1474 12529 1502 13667
rect 2338 13149 2366 13713
rect 2338 13121 2462 13149
rect 2434 12973 2462 13121
rect 2626 12927 2654 14157
rect 2434 12899 2654 12927
rect 1282 12455 1406 12483
rect 1378 12307 1406 12455
rect 994 12233 1214 12261
rect 1186 11641 1214 12233
rect 2434 12187 2462 12899
rect 2434 12159 2558 12187
rect 1378 11197 1406 11743
rect 34 10753 158 10781
rect 34 9523 62 10753
rect 1090 10531 1118 10781
rect 994 10115 1022 10263
rect 898 10087 1022 10115
rect 0 9495 97 9523
rect 898 9227 926 10087
rect 898 9199 1022 9227
rect 994 9051 1022 9199
rect 34 8977 158 9005
rect 34 8117 62 8977
rect 1186 8533 1214 10337
rect 1474 9523 1502 10337
rect 1378 9495 1502 9523
rect 1378 8755 1406 9495
rect 1474 8977 1502 9449
rect 1858 9199 1886 9597
rect 0 8089 97 8117
rect 706 7201 734 7747
rect 1090 7201 1118 8265
rect 1858 7867 1886 8191
rect 1954 7821 1982 11447
rect 2050 9199 2078 9597
rect 2242 8413 2270 12113
rect 2530 10929 2558 12159
rect 2434 10901 2558 10929
rect 2434 10309 2462 10901
rect 3202 10235 3230 14925
rect 2434 9643 2462 10115
rect 3106 8977 3134 10115
rect 3298 9199 3326 9449
rect 2914 8857 2942 8931
rect 3490 8857 3518 15119
rect 4258 13565 4286 14851
rect 4354 14703 4382 17663
rect 4546 17191 4574 22103
rect 4834 20475 4862 22149
rect 5410 21187 5438 21659
rect 5794 20845 5822 22177
rect 5986 21631 6014 23407
rect 6274 22519 6302 26173
rect 7810 26099 7838 27181
rect 7906 27033 8030 27061
rect 7906 26293 7934 27033
rect 6466 25627 6494 26099
rect 7810 26071 7934 26099
rect 6658 24295 6686 25729
rect 7906 24443 7934 26071
rect 8098 25849 8126 26987
rect 8290 26885 8318 27653
rect 8578 27061 8606 27699
rect 8482 27033 8606 27061
rect 9154 27061 9182 27773
rect 9154 27033 9278 27061
rect 8290 26367 8318 26765
rect 8482 25877 8510 27033
rect 8386 25849 8510 25877
rect 8098 24517 8126 25063
rect 8386 24961 8414 25849
rect 8674 25137 8702 26913
rect 9250 26885 9278 27033
rect 9442 26765 9470 28319
rect 9346 26737 9470 26765
rect 9346 26025 9374 26737
rect 9346 25997 9470 26025
rect 9442 25849 9470 25997
rect 9634 25729 9662 28439
rect 9826 28171 9854 28985
rect 9826 28143 9950 28171
rect 9922 27579 9950 28143
rect 9826 27551 9950 27579
rect 9826 27181 9854 27551
rect 9826 26765 9854 26913
rect 9826 26737 9950 26765
rect 9922 26173 9950 26737
rect 9538 25701 9662 25729
rect 9826 26145 9950 26173
rect 8674 25109 8798 25137
rect 8290 24397 8318 24767
rect 8194 24369 8318 24397
rect 6946 24175 6974 24323
rect 6658 24147 6782 24175
rect 6946 24147 7070 24175
rect 6082 21853 6110 22399
rect 5794 20817 5918 20845
rect 4738 20447 4862 20475
rect 4738 20299 4766 20447
rect 4738 17635 4766 19809
rect 4930 19143 4958 20105
rect 5602 19633 5630 20771
rect 5890 20253 5918 20817
rect 5794 20225 5918 20253
rect 6274 20225 6302 21881
rect 6754 21705 6782 24147
rect 7042 23657 7070 24147
rect 6946 23629 7070 23657
rect 6946 23185 6974 23629
rect 7138 21631 7166 23509
rect 7906 22297 7934 24101
rect 8194 23879 8222 24369
rect 8194 23851 8318 23879
rect 8290 23703 8318 23851
rect 8482 23435 8510 25063
rect 8770 24323 8798 25109
rect 9538 24915 9566 25701
rect 9538 24887 9662 24915
rect 8674 24295 8798 24323
rect 9442 24295 9470 24767
rect 8674 24147 8702 24295
rect 8386 23407 8510 23435
rect 8386 22473 8414 23407
rect 8770 23361 8798 23731
rect 8674 23333 8798 23361
rect 8674 22519 8702 23333
rect 9058 23037 9086 24175
rect 8386 22445 8510 22473
rect 8098 21853 8126 22251
rect 6562 20373 6590 20771
rect 5794 19735 5822 20225
rect 5794 19707 5918 19735
rect 4930 19115 5054 19143
rect 5026 18181 5054 19115
rect 5794 19069 5822 19217
rect 4930 18153 5054 18181
rect 5698 19041 5822 19069
rect 4930 17635 4958 18153
rect 5698 17737 5726 19041
rect 5986 17783 6014 20105
rect 6178 19439 6206 19587
rect 6754 19559 6782 21585
rect 6946 20965 6974 21437
rect 7330 21187 7358 21659
rect 6946 19707 6974 20845
rect 7138 19855 7166 20919
rect 7330 19735 7358 20993
rect 8290 20521 8318 20771
rect 7522 20179 7550 20327
rect 7522 20151 7646 20179
rect 7234 19707 7358 19735
rect 6178 19411 6302 19439
rect 6274 18847 6302 19411
rect 6178 18819 6302 18847
rect 6178 18301 6206 18819
rect 7234 18699 7262 19707
rect 7618 19661 7646 20151
rect 7522 19633 7646 19661
rect 7522 18773 7550 19633
rect 7522 18745 7646 18773
rect 7234 18671 7358 18699
rect 7330 18523 7358 18671
rect 5698 17709 5822 17737
rect 4642 16303 4670 16923
rect 4834 16525 4862 16997
rect 5794 16895 5822 17709
rect 7330 17635 7358 18329
rect 7618 18181 7646 18745
rect 7522 18153 7646 18181
rect 7522 17811 7550 18153
rect 7522 17783 7646 17811
rect 6178 17561 6302 17589
rect 4354 14675 4574 14703
rect 4546 13565 4574 14675
rect 5122 14453 5150 15665
rect 5602 14527 5630 15665
rect 6082 14527 6110 14925
rect 5410 14083 5438 14407
rect 6274 14231 6302 17561
rect 6658 16895 6686 17515
rect 7330 17117 7358 17515
rect 7618 17071 7646 17783
rect 7906 17191 7934 18773
rect 8098 18449 8126 19735
rect 8482 18403 8510 22445
rect 9250 22399 9278 23583
rect 9154 22371 9278 22399
rect 9154 21659 9182 22371
rect 9442 21705 9470 23657
rect 9154 21631 9278 21659
rect 8674 20845 8702 20993
rect 8674 20817 8798 20845
rect 8770 20327 8798 20817
rect 9058 20521 9086 20771
rect 8674 20299 8798 20327
rect 8674 20151 8702 20299
rect 8962 19513 8990 19661
rect 8866 19485 8990 19513
rect 8866 18921 8894 19485
rect 9058 18967 9086 20253
rect 8866 18893 8990 18921
rect 8962 18773 8990 18893
rect 8962 18745 9086 18773
rect 8482 18375 8990 18403
rect 7522 17043 7646 17071
rect 6850 14379 6878 15443
rect 5506 13639 5534 14111
rect 7042 13861 7070 14407
rect 7234 14185 7262 16331
rect 7522 14379 7550 17043
rect 7810 15563 7838 16405
rect 8098 16377 8126 16775
rect 8386 16525 8414 16997
rect 8482 16155 8510 18255
rect 8962 17635 8990 18375
rect 9058 18301 9086 18745
rect 8674 17145 8702 17441
rect 8674 17117 8798 17145
rect 8770 16553 8798 17117
rect 8674 16525 8798 16553
rect 9058 16525 9086 16849
rect 8674 16377 8702 16525
rect 9250 16229 9278 21631
rect 9634 20965 9662 24887
rect 9826 23139 9854 26145
rect 10306 25849 10334 26099
rect 10690 25729 10718 25877
rect 10594 25701 10718 25729
rect 10594 25137 10622 25701
rect 10594 25109 10718 25137
rect 10114 23851 10142 24249
rect 10594 24221 10622 24989
rect 10690 24961 10718 25109
rect 10882 24101 10910 26913
rect 11458 26469 11486 29059
rect 11650 28911 11678 29623
rect 11938 29179 11966 29577
rect 11650 28883 11870 28911
rect 11842 28615 11870 28883
rect 11746 28587 11870 28615
rect 11746 27801 11774 28587
rect 12034 27847 12062 28911
rect 11746 27773 11870 27801
rect 11842 26959 11870 27773
rect 12610 27431 12638 28097
rect 13474 27579 13502 31575
rect 13954 29031 13982 30095
rect 13858 28735 13982 28763
rect 13474 27551 13790 27579
rect 12610 27403 12734 27431
rect 11362 26441 11486 26469
rect 11362 25803 11390 26441
rect 11362 25775 11486 25803
rect 11458 25627 11486 25775
rect 9826 23111 9950 23139
rect 9922 22547 9950 23111
rect 9826 22519 9950 22547
rect 9826 22371 9854 22519
rect 9826 21807 9854 22251
rect 9826 21779 9950 21807
rect 9922 20919 9950 21779
rect 10306 21631 10334 24101
rect 10786 24073 10910 24101
rect 10786 23509 10814 24073
rect 11074 23555 11102 25433
rect 11458 23805 11486 24915
rect 11650 24887 11678 26913
rect 11362 23777 11486 23805
rect 10786 23481 10910 23509
rect 9826 20891 9950 20919
rect 9538 20299 9566 20771
rect 9538 19365 9566 19513
rect 9442 19337 9566 19365
rect 9442 18551 9470 19337
rect 9442 18523 9566 18551
rect 9538 18375 9566 18523
rect 9634 17487 9662 20253
rect 9826 19143 9854 20891
rect 10018 20327 10046 20475
rect 10018 20299 10142 20327
rect 10114 19809 10142 20299
rect 10498 19855 10526 21659
rect 10882 21631 10910 23481
rect 11362 22843 11390 23777
rect 11362 22815 11486 22843
rect 11458 22297 11486 22815
rect 11458 20965 11486 21659
rect 11458 20373 11486 20771
rect 11650 19809 11678 24175
rect 12034 23851 12062 24989
rect 12226 24961 12254 26247
rect 12706 26219 12734 27403
rect 13282 27283 13310 27431
rect 13186 27255 13310 27283
rect 13186 26543 13214 27255
rect 13186 26515 13310 26543
rect 12994 24295 13022 25729
rect 13282 24175 13310 26515
rect 13474 26469 13502 27551
rect 13858 26515 13886 28735
rect 14050 27847 14078 28245
rect 14530 27505 14558 29651
rect 16258 28735 16286 29429
rect 16450 29105 16478 29651
rect 16642 28883 16670 29577
rect 17026 27625 17054 30317
rect 17122 29845 17150 30317
rect 18658 27699 18686 28245
rect 14434 27477 14558 27505
rect 13474 26441 13598 26469
rect 13570 25877 13598 26441
rect 13474 25849 13598 25877
rect 13474 25137 13502 25849
rect 14434 25803 14462 27477
rect 14434 25775 14558 25803
rect 14530 25433 14558 25775
rect 14722 25729 14750 27431
rect 16738 26515 16766 27505
rect 20674 26515 20702 28319
rect 21154 27801 21182 28097
rect 21154 27773 21278 27801
rect 20962 26885 20990 27727
rect 21250 26839 21278 27773
rect 21154 26811 21278 26839
rect 14722 25701 14846 25729
rect 13474 25109 13598 25137
rect 13570 24175 13598 25109
rect 13186 24147 13310 24175
rect 13474 24147 13598 24175
rect 11842 23287 11870 23435
rect 11842 23259 11966 23287
rect 11938 22547 11966 23259
rect 11842 22519 11966 22547
rect 11842 22371 11870 22519
rect 12706 22325 12734 23657
rect 13186 23509 13214 24147
rect 12610 22297 12734 22325
rect 12706 21733 12734 22297
rect 12610 21705 12734 21733
rect 12994 23481 13214 23509
rect 11842 21187 11870 21437
rect 12034 20919 12062 21659
rect 11986 20891 12062 20919
rect 12610 20919 12638 21705
rect 12802 21631 12926 21659
rect 12898 20965 12926 21631
rect 12994 21039 13022 23481
rect 13282 23185 13310 23435
rect 12610 20891 12734 20919
rect 10018 19781 10142 19809
rect 11554 19781 11678 19809
rect 10018 19633 10046 19781
rect 11554 19217 11582 19781
rect 11554 19189 11678 19217
rect 11842 19189 11870 20475
rect 11986 20327 12014 20891
rect 12130 20373 12158 20771
rect 11986 20299 12062 20327
rect 9826 19115 9950 19143
rect 9922 18477 9950 19115
rect 11650 19069 11678 19189
rect 12034 19115 12062 20299
rect 12706 19781 12734 20891
rect 11650 19041 11774 19069
rect 9826 18449 9950 18477
rect 9826 17857 9854 18449
rect 11458 18227 11486 18995
rect 11746 18181 11774 19041
rect 11650 18153 11774 18181
rect 12034 18967 12158 18995
rect 10402 17635 10430 18107
rect 11650 17663 11678 18153
rect 11650 17635 11774 17663
rect 9442 16997 9470 17145
rect 9442 16969 9566 16997
rect 9538 16479 9566 16969
rect 10114 16775 10142 17589
rect 9442 16451 9566 16479
rect 9442 16303 9470 16451
rect 9250 15711 9278 16109
rect 9826 15859 9854 16775
rect 10114 16747 10334 16775
rect 10786 16747 10814 17589
rect 11650 17191 11678 17635
rect 12034 17117 12062 18967
rect 12130 16895 12158 17663
rect 12322 17145 12350 19735
rect 12706 19189 12734 19513
rect 13090 18995 13118 21659
rect 13474 20373 13502 24147
rect 13858 21409 13886 22991
rect 14146 21853 14174 24767
rect 14338 24443 14366 24915
rect 14434 24517 14462 25433
rect 14530 25405 14654 25433
rect 14338 21853 14366 22769
rect 14626 22371 14654 25405
rect 14914 25183 14942 25655
rect 16162 25405 16190 26099
rect 15202 23185 15230 23583
rect 15490 23185 15518 24323
rect 15682 23629 15710 25063
rect 16450 23703 16478 26321
rect 18466 25627 18494 26321
rect 16642 22917 16670 23065
rect 16546 22889 16670 22917
rect 16546 22399 16574 22889
rect 16546 22371 16670 22399
rect 14626 20151 14654 20993
rect 15202 20225 15230 22103
rect 16642 21733 16670 22371
rect 16450 21705 16670 21733
rect 16834 21733 16862 24767
rect 18946 24323 18974 25655
rect 19426 25627 19454 26099
rect 19906 25849 19934 26321
rect 20194 25183 20222 25729
rect 19138 24767 19166 24915
rect 19138 24739 19262 24767
rect 18850 24295 18974 24323
rect 17794 23037 17822 23435
rect 18850 23139 18878 24295
rect 19234 24249 19262 24739
rect 20386 24369 20414 25729
rect 21154 24369 21182 26811
rect 21634 26765 21662 26913
rect 21538 26737 21662 26765
rect 21538 26025 21566 26737
rect 21538 25997 21662 26025
rect 21634 25849 21662 25997
rect 21634 24841 21662 24989
rect 21538 24813 21662 24841
rect 21538 24323 21566 24813
rect 19138 24221 19262 24249
rect 18850 23111 18974 23139
rect 17506 22445 17534 22991
rect 18946 22843 18974 23111
rect 18850 22815 18974 22843
rect 17122 21853 17150 22325
rect 18850 21779 18878 22815
rect 19138 22251 19166 24221
rect 19906 22519 19934 24323
rect 21538 24295 21662 24323
rect 20194 22889 20222 24101
rect 21634 24027 21662 24295
rect 21538 23999 21662 24027
rect 21538 23065 21566 23999
rect 21826 23139 21854 31057
rect 22306 26839 22334 29503
rect 24034 28171 24062 28467
rect 24034 28143 24158 28171
rect 23746 27283 23774 27431
rect 22210 26811 22334 26839
rect 23650 27255 23774 27283
rect 22210 26173 22238 26811
rect 22498 26247 22526 26765
rect 23650 26691 23678 27255
rect 23650 26663 23774 26691
rect 23746 26515 23774 26663
rect 22498 26219 22622 26247
rect 22210 26145 22334 26173
rect 22306 25803 22334 26145
rect 22210 25775 22334 25803
rect 22210 24915 22238 25775
rect 22594 25729 22622 26219
rect 22498 25701 22622 25729
rect 23170 25701 23198 26247
rect 23938 26145 23966 27431
rect 24130 27135 24158 28143
rect 24130 27107 24254 27135
rect 24226 26173 24254 27107
rect 24130 26145 24254 26173
rect 22498 24961 22526 25701
rect 22210 24887 22334 24915
rect 21826 23111 21950 23139
rect 21538 23037 21662 23065
rect 21250 22371 21278 22769
rect 21442 22251 21470 22917
rect 19042 22223 19166 22251
rect 21346 22223 21470 22251
rect 16834 21705 16958 21733
rect 16450 21141 16478 21705
rect 16354 21113 16478 21141
rect 16354 20179 16382 21113
rect 16354 20151 16478 20179
rect 14050 20077 14174 20105
rect 12514 18523 12542 18995
rect 13090 18967 13310 18995
rect 13090 18819 13214 18847
rect 12706 17191 12734 17515
rect 12322 17117 12542 17145
rect 10306 16525 10334 16747
rect 12322 16303 12350 17117
rect 12706 16377 12734 16775
rect 7234 14157 7454 14185
rect 7234 13741 7262 14111
rect 7138 13713 7262 13741
rect 3682 12899 3710 13445
rect 7138 13075 7166 13713
rect 2722 8829 2942 8857
rect 3394 8829 3518 8857
rect 2242 8385 2366 8413
rect 1858 7793 1982 7821
rect 1858 7007 1886 7793
rect 2146 7201 2174 8339
rect 226 6785 254 6859
rect 0 6757 254 6785
rect 706 5869 734 6933
rect 34 5647 158 5675
rect 34 5453 62 5647
rect 1474 5573 1502 6859
rect 1762 6785 1790 7007
rect 1858 6979 1982 7007
rect 1762 6757 1886 6785
rect 0 5425 97 5453
rect 34 4315 158 4343
rect 34 4121 62 4315
rect 0 4093 97 4121
rect 1474 3751 1502 5453
rect 1858 4537 1886 6757
rect 1954 6387 1982 6979
rect 2146 5203 2174 6785
rect 2338 6535 2366 8385
rect 2722 8311 2750 8829
rect 3394 8265 3422 8829
rect 2338 4981 2366 5601
rect 2626 5129 2654 8265
rect 3394 8237 3518 8265
rect 3298 7719 3326 8117
rect 3490 7599 3518 8237
rect 3394 7571 3518 7599
rect 2722 4537 2750 5601
rect 3106 5573 3134 7451
rect 3394 6711 3422 7571
rect 3394 6683 3518 6711
rect 3490 6535 3518 6683
rect 3298 6267 3326 6415
rect 3298 6239 3422 6267
rect 3394 5749 3422 6239
rect 3298 5721 3422 5749
rect 3298 5601 3326 5721
rect 3202 5573 3326 5601
rect 3202 5453 3230 5573
rect 3010 5425 3230 5453
rect 3010 4861 3038 5425
rect 3010 4833 3134 4861
rect 1474 3723 1598 3751
rect 2434 3649 2462 4269
rect 34 3501 158 3529
rect 34 2715 62 3501
rect 2818 3455 2846 4417
rect 3106 4389 3134 4833
rect 3010 3871 3038 4343
rect 2818 3427 3134 3455
rect 3106 2983 3134 3427
rect 3298 3205 3326 5083
rect 0 2687 97 2715
rect 34 1383 62 1679
rect 2722 1651 2750 2271
rect 3106 1873 3134 2419
rect 3394 1651 3422 2345
rect 3490 2169 3518 4343
rect 3682 3825 3710 10781
rect 3874 9865 3902 12261
rect 4354 10411 4382 10929
rect 4258 10383 4382 10411
rect 3778 8533 3806 9671
rect 4258 9523 4286 10383
rect 4258 9495 4382 9523
rect 4162 8857 4190 9005
rect 4066 8829 4190 8857
rect 4066 8265 4094 8829
rect 4354 8459 4382 9495
rect 4546 9199 4574 10337
rect 4642 10263 4670 11447
rect 4834 10309 4862 12779
rect 5026 12187 5054 12335
rect 5026 12159 5150 12187
rect 5122 11521 5150 12159
rect 5026 11493 5150 11521
rect 5026 11151 5054 11493
rect 5026 11123 5150 11151
rect 5122 10485 5150 11123
rect 5026 10457 5150 10485
rect 5026 10337 5054 10457
rect 4930 10309 5054 10337
rect 4642 10235 4766 10263
rect 4066 8237 4190 8265
rect 4162 8117 4190 8237
rect 4162 8089 4286 8117
rect 4258 7895 4286 8089
rect 4066 7867 4286 7895
rect 4066 7053 4094 7867
rect 4354 7821 4382 8339
rect 4258 7793 4382 7821
rect 3970 5647 3998 6267
rect 4258 5721 4286 7793
rect 4546 6461 4574 9005
rect 4738 6387 4766 10235
rect 4930 9717 4958 10309
rect 5122 9199 5150 10337
rect 5506 9819 5534 12779
rect 5794 12529 5822 13075
rect 7138 13047 7262 13075
rect 7234 12927 7262 13047
rect 5794 10189 5822 11743
rect 5410 9791 5534 9819
rect 5698 10161 5822 10189
rect 5410 9301 5438 9791
rect 5698 9375 5726 10161
rect 5698 9347 5822 9375
rect 5410 9273 5534 9301
rect 4834 8829 4862 9005
rect 4930 7719 4958 8339
rect 5122 7201 5150 8265
rect 5506 7747 5534 9273
rect 5794 9199 5822 9347
rect 5506 7719 5726 7747
rect 5506 7201 5534 7673
rect 5698 7155 5726 7719
rect 5602 7127 5726 7155
rect 4930 6535 4958 7007
rect 5026 6489 5054 6785
rect 4930 6461 5054 6489
rect 4930 5869 4958 6461
rect 5602 5749 5630 7127
rect 5506 5721 5630 5749
rect 5890 5749 5918 10115
rect 5890 5721 6014 5749
rect 3874 5203 3902 5453
rect 5506 5083 5534 5721
rect 5794 5129 5822 5675
rect 5986 5083 6014 5721
rect 3682 3797 3806 3825
rect 3778 2863 3806 3797
rect 4642 3723 4670 4121
rect 3682 2835 3806 2863
rect 0 1355 97 1383
rect 3682 1235 3710 2835
rect 4546 1725 4574 3529
rect 3586 1207 3710 1235
rect 4834 1207 4862 5083
rect 5506 5055 5630 5083
rect 5122 3871 5150 5009
rect 5602 2493 5630 5055
rect 5890 5055 6014 5083
rect 5890 2539 5918 5055
rect 6178 3649 6206 12113
rect 6850 11521 6878 12187
rect 7138 11863 7166 12927
rect 7234 12899 7310 12927
rect 7282 11891 7310 12899
rect 7426 12483 7454 14157
rect 7426 12455 7550 12483
rect 7234 11863 7310 11891
rect 7234 11743 7262 11863
rect 6754 11493 6878 11521
rect 6754 10855 6782 11493
rect 6754 10827 6878 10855
rect 6850 10383 6878 10827
rect 6466 8117 6494 9153
rect 6658 8533 6686 9005
rect 6850 8339 6878 9449
rect 6850 8311 6974 8339
rect 6466 8089 6686 8117
rect 6370 5869 6398 6341
rect 6658 5795 6686 8089
rect 6850 7645 6878 8311
rect 7042 7719 7070 11743
rect 7234 11715 7358 11743
rect 7234 10337 7262 11715
rect 7522 11521 7550 12455
rect 7906 12261 7934 14925
rect 7906 12233 8030 12261
rect 7906 12113 7934 12233
rect 7426 11493 7550 11521
rect 7810 12085 7934 12113
rect 7810 11521 7838 12085
rect 7810 11493 7934 11521
rect 7426 11151 7454 11493
rect 7426 11123 7550 11151
rect 7138 10309 7262 10337
rect 7522 10189 7550 11123
rect 7906 10411 7934 11493
rect 8098 11197 8126 14111
rect 8290 12187 8318 15591
rect 10978 14527 11006 16257
rect 13090 15785 13118 18819
rect 13282 18523 13310 18967
rect 13474 17635 13502 19439
rect 14050 19365 14078 20077
rect 13954 19337 14078 19365
rect 13954 18847 13982 19337
rect 14242 19069 14270 19439
rect 14242 19041 14366 19069
rect 13954 18819 14078 18847
rect 14050 18477 14078 18819
rect 13954 18449 14078 18477
rect 13954 17737 13982 18449
rect 13954 17709 14078 17737
rect 14050 17561 14078 17709
rect 14242 17561 14270 19041
rect 14626 18995 14654 19661
rect 16450 19559 16478 20151
rect 16642 20077 16670 21659
rect 16930 20401 16958 21705
rect 17506 20521 17534 20993
rect 16834 20373 16958 20401
rect 16834 20225 16862 20373
rect 18178 20225 18206 21585
rect 19042 20373 19070 22223
rect 19618 20891 19646 21585
rect 20098 20521 20126 21659
rect 20290 21187 20318 21659
rect 17026 19189 17054 19661
rect 14626 18967 14846 18995
rect 14626 18375 14654 18967
rect 16258 18523 16286 18995
rect 16930 18181 16958 19069
rect 17410 18523 17438 18773
rect 16834 18153 16958 18181
rect 12130 15443 12158 15591
rect 11938 15415 12158 15443
rect 11938 14703 11966 15415
rect 12226 15147 12254 15443
rect 12226 15119 12446 15147
rect 11938 14675 12158 14703
rect 12130 14527 12158 14675
rect 9634 13713 9662 14111
rect 10306 13741 10334 14333
rect 10114 13713 10334 13741
rect 10114 12853 10142 13713
rect 10114 12825 10334 12853
rect 10402 12825 10430 13667
rect 10594 13519 10622 14259
rect 10546 13491 10622 13519
rect 10546 13001 10574 13491
rect 10690 13047 10718 13445
rect 11458 13195 11486 13667
rect 11554 13565 11582 14259
rect 12034 13787 12062 14333
rect 12418 14259 12446 15119
rect 12706 14527 12734 14999
rect 12994 14971 13022 15665
rect 13186 15119 13214 15591
rect 14050 14851 14078 16183
rect 15106 15637 15134 17145
rect 15202 17043 15230 17441
rect 15394 17043 15422 17441
rect 15490 16303 15518 17589
rect 15682 16183 15710 17737
rect 16834 17589 16862 18153
rect 16834 17561 16958 17589
rect 17026 17561 17054 18107
rect 17506 17635 17534 18329
rect 16930 17413 16958 17561
rect 17890 17117 17918 18921
rect 15586 16155 15710 16183
rect 15586 15369 15614 16155
rect 15586 15341 15710 15369
rect 15682 15073 15710 15341
rect 13954 14823 14078 14851
rect 15586 15045 15710 15073
rect 13954 14407 13982 14823
rect 13858 14379 13982 14407
rect 12226 14231 12446 14259
rect 12226 13593 12254 14231
rect 11746 13565 12254 13593
rect 10546 12973 10622 13001
rect 9730 12307 9758 12779
rect 10306 12381 10334 12825
rect 8290 12159 8414 12187
rect 8386 11151 8414 12159
rect 8290 11123 8414 11151
rect 7906 10383 8222 10411
rect 7330 10161 7550 10189
rect 7330 9153 7358 10161
rect 8194 9643 8222 10383
rect 8290 10337 8318 11123
rect 8674 10383 8702 11447
rect 8866 11197 8894 11669
rect 8290 10309 8414 10337
rect 7618 9199 7646 9597
rect 8002 9199 8030 9597
rect 7330 9125 7934 9153
rect 7234 8857 7262 9005
rect 7234 8829 7358 8857
rect 7330 8043 7358 8829
rect 7234 8015 7358 8043
rect 7042 7007 7070 7155
rect 6946 6979 7070 7007
rect 7234 7007 7262 8015
rect 7234 6979 7358 7007
rect 6946 6489 6974 6979
rect 7234 6535 7262 6785
rect 6946 6461 7070 6489
rect 6658 3205 6686 5083
rect 7042 4907 7070 6461
rect 7906 6341 7934 9125
rect 8194 6979 8222 8339
rect 8386 7599 8414 10309
rect 9058 9523 9086 11743
rect 9634 9745 9662 12187
rect 10402 11863 10430 12261
rect 10594 11641 10622 12973
rect 10882 11521 10910 12483
rect 10786 11493 10910 11521
rect 9922 10531 9950 10781
rect 10786 10485 10814 11493
rect 10786 10457 10910 10485
rect 10882 10309 10910 10457
rect 9634 9717 9758 9745
rect 9058 9495 9182 9523
rect 8962 8265 8990 8857
rect 9058 8311 9086 9449
rect 9154 9051 9182 9495
rect 8962 8237 9086 8265
rect 8674 7719 8702 8117
rect 9058 7821 9086 8237
rect 9442 8191 9470 9671
rect 9730 9079 9758 9717
rect 9634 9051 9758 9079
rect 10594 9051 10622 10115
rect 11074 9227 11102 12261
rect 11554 11669 11582 11817
rect 11458 11641 11582 11669
rect 11458 10929 11486 11641
rect 11458 10901 11582 10929
rect 11746 10901 11774 13565
rect 12994 13195 13022 14333
rect 13186 13861 13214 14333
rect 13858 13001 13886 14379
rect 12034 12085 12158 12113
rect 12034 10901 12062 12085
rect 11458 9643 11486 10781
rect 11554 10531 11582 10901
rect 12322 10383 12350 12409
rect 12706 12261 12734 13001
rect 13762 12973 13886 13001
rect 12706 12233 12830 12261
rect 12706 12113 12734 12233
rect 12610 12085 12734 12113
rect 12610 11521 12638 12085
rect 12610 11493 12734 11521
rect 12706 10235 12734 11493
rect 12898 11197 12926 12335
rect 13186 11567 13214 12557
rect 13762 12261 13790 12973
rect 14146 12927 14174 14777
rect 15586 14481 15614 15045
rect 15586 14453 15710 14481
rect 14530 13195 14558 14333
rect 15682 14305 15710 14453
rect 14050 12899 14174 12927
rect 13762 12233 13886 12261
rect 13858 12085 13886 12233
rect 12994 10531 13022 10929
rect 13186 10411 13214 11447
rect 13762 10975 13790 11817
rect 14050 11197 14078 12899
rect 13090 10383 13214 10411
rect 11746 9643 11774 10115
rect 13090 9745 13118 10383
rect 13090 9717 13214 9745
rect 11074 9199 11198 9227
rect 9634 8903 9662 9051
rect 10306 8459 10334 9005
rect 9442 8163 9566 8191
rect 8962 7793 9086 7821
rect 8386 7571 8510 7599
rect 8194 6637 8222 6785
rect 8194 6609 8270 6637
rect 7906 6313 8126 6341
rect 6946 3723 6974 4787
rect 7906 3899 7934 6267
rect 8098 5675 8126 6313
rect 8242 5897 8270 6609
rect 8482 6563 8510 7571
rect 8962 6859 8990 7793
rect 9250 6859 9278 8117
rect 9538 7377 9566 8163
rect 10978 7867 11006 9005
rect 11554 8977 11582 9523
rect 12802 9449 12830 9597
rect 12706 9421 12830 9449
rect 11650 7793 11678 9005
rect 9442 7349 9566 7377
rect 9442 7201 9470 7349
rect 9730 6859 9758 7007
rect 8962 6831 9086 6859
rect 9250 6831 9374 6859
rect 8386 6535 8510 6563
rect 8386 6239 8414 6535
rect 8194 5869 8270 5897
rect 8194 5721 8222 5869
rect 8098 5647 8222 5675
rect 7810 3871 7934 3899
rect 7810 3649 7838 3871
rect 8194 3751 8222 5647
rect 8578 4315 8606 5453
rect 8674 5203 8702 6415
rect 9058 6045 9086 6831
rect 9346 6267 9374 6831
rect 9250 6239 9374 6267
rect 9634 6831 9758 6859
rect 9922 6933 9950 7673
rect 10402 7201 10430 7451
rect 11746 7201 11774 7747
rect 11938 7645 11966 8931
rect 12130 8459 12158 9079
rect 12706 8857 12734 9421
rect 12706 8829 12830 8857
rect 12802 8533 12830 8829
rect 12130 8043 12158 8339
rect 12034 8015 12158 8043
rect 12034 7599 12062 8015
rect 12994 7867 13022 9597
rect 13186 8533 13214 9717
rect 13378 9153 13406 10855
rect 14242 10383 14270 11669
rect 13954 9199 13982 10263
rect 14530 10161 14558 12779
rect 15106 12455 15134 12927
rect 15298 12557 15326 14111
rect 15874 13565 15902 16775
rect 16258 14379 16286 16109
rect 16930 15637 16958 16997
rect 18178 16525 18206 16997
rect 18754 16895 18782 19587
rect 18658 16553 18686 16775
rect 18658 16525 18782 16553
rect 17122 15711 17150 16331
rect 17410 15711 17438 16183
rect 17794 15859 17822 16257
rect 18274 15859 18302 16331
rect 16546 15517 16574 15591
rect 16450 15489 16574 15517
rect 16450 13639 16478 15489
rect 17506 15147 17534 15739
rect 18658 15637 18686 16331
rect 18754 15591 18782 16525
rect 18658 15563 18782 15591
rect 17410 15119 17534 15147
rect 17410 14185 17438 15119
rect 17698 14407 17726 15147
rect 17650 14379 17726 14407
rect 17410 14157 17534 14185
rect 17506 13787 17534 14157
rect 17650 13667 17678 14379
rect 17794 13861 17822 14333
rect 17602 13639 17678 13667
rect 16258 13149 16286 13445
rect 16162 13121 16286 13149
rect 15298 12529 15422 12557
rect 14818 12039 14846 12335
rect 16162 12187 16190 13121
rect 17602 13075 17630 13639
rect 17890 13121 17918 13667
rect 18082 13565 18110 14407
rect 18658 14157 18686 15563
rect 19042 15443 19070 17441
rect 18946 15415 19070 15443
rect 18946 14703 18974 15415
rect 19234 15295 19262 15443
rect 19186 15267 19262 15295
rect 18946 14675 19070 14703
rect 19042 14527 19070 14675
rect 19186 14407 19214 15267
rect 19330 14453 19358 17811
rect 19522 16479 19550 20253
rect 19810 16775 19838 17663
rect 19906 17635 19934 18107
rect 19810 16747 19934 16775
rect 19522 16451 19646 16479
rect 19618 15517 19646 16451
rect 19906 16229 19934 16747
rect 20098 16525 20126 18255
rect 19522 15489 19646 15517
rect 19522 15147 19550 15489
rect 19522 15119 19646 15147
rect 19618 14407 19646 15119
rect 19186 14379 19262 14407
rect 18274 13223 18302 14111
rect 19042 13565 19070 14111
rect 19234 13741 19262 14379
rect 19186 13713 19262 13741
rect 19522 14379 19646 14407
rect 19522 13741 19550 14379
rect 19522 13713 19646 13741
rect 18274 13195 18494 13223
rect 16162 12159 16286 12187
rect 14722 12011 14846 12039
rect 14722 10901 14750 12011
rect 16258 11817 16286 12159
rect 16162 11789 16286 11817
rect 15490 11077 15518 11595
rect 16162 11077 16190 11789
rect 16450 11151 16478 13075
rect 17602 13047 17726 13075
rect 16546 12455 16574 13001
rect 16930 11715 16958 12779
rect 17698 12039 17726 13047
rect 17602 12011 17726 12039
rect 17602 11521 17630 12011
rect 17986 11965 18014 12113
rect 17890 11937 18014 11965
rect 17602 11493 17726 11521
rect 16450 11123 16574 11151
rect 17698 11123 17726 11493
rect 15490 11049 15614 11077
rect 16162 11049 16286 11077
rect 13378 9125 13502 9153
rect 13474 8487 13502 9125
rect 15298 9051 15326 11003
rect 15586 10485 15614 11049
rect 16258 10901 16286 11049
rect 15490 10457 15614 10485
rect 15490 10309 15518 10457
rect 16258 10263 16286 10781
rect 16162 10235 16286 10263
rect 16162 9523 16190 10235
rect 16546 10189 16574 11123
rect 17698 10531 17726 10929
rect 17890 10855 17918 11937
rect 18082 10901 18110 12335
rect 18274 11817 18302 12853
rect 18466 12529 18494 13195
rect 18850 13047 18878 13445
rect 19042 12307 19070 13445
rect 19186 12187 19214 13713
rect 19330 13149 19358 13667
rect 19330 13121 19454 13149
rect 19330 12233 19358 13121
rect 19618 12853 19646 13713
rect 19906 13639 19934 15591
rect 20098 13713 20126 15887
rect 20290 15443 20318 18921
rect 20386 18893 20414 21585
rect 21346 21215 21374 22223
rect 21346 21187 21470 21215
rect 21442 21039 21470 21187
rect 21634 20919 21662 23037
rect 21922 22177 21950 23111
rect 21826 22149 21950 22177
rect 21826 21807 21854 22149
rect 21826 21779 21950 21807
rect 21538 20891 21662 20919
rect 21250 19041 21278 20327
rect 21538 18477 21566 20891
rect 21922 20845 21950 21779
rect 22306 21631 22334 24887
rect 22594 23185 22622 24323
rect 22594 21187 22622 22547
rect 22978 22519 23006 22917
rect 23074 20891 23102 22325
rect 23458 20965 23486 24397
rect 23650 24369 23678 25729
rect 24130 24175 24158 26145
rect 24034 24147 24158 24175
rect 24034 23139 24062 24147
rect 24034 23111 24158 23139
rect 24130 22963 24158 23111
rect 24034 22325 24062 22917
rect 24226 22843 24254 22991
rect 23938 22297 24062 22325
rect 24178 22815 24254 22843
rect 24178 22325 24206 22815
rect 24322 22371 24350 24101
rect 24178 22297 24254 22325
rect 23938 21807 23966 22297
rect 23938 21779 24062 21807
rect 24226 21779 24254 22297
rect 24034 21631 24062 21779
rect 21826 20817 21950 20845
rect 21538 18449 21662 18477
rect 21634 18301 21662 18449
rect 20482 16895 20510 18107
rect 21826 17663 21854 20817
rect 22402 19189 22430 20253
rect 23074 19707 23102 20771
rect 23650 19217 23678 21067
rect 24130 20919 24158 21437
rect 23650 19189 23774 19217
rect 22114 18227 22142 19069
rect 23746 17709 23774 19189
rect 21826 17635 21950 17663
rect 20578 15563 20606 16849
rect 21058 16257 21086 17441
rect 21442 16701 21470 17441
rect 21634 16997 21662 17589
rect 20962 16229 21086 16257
rect 21346 16673 21470 16701
rect 21538 16969 21662 16997
rect 21346 16109 21374 16673
rect 21250 16081 21374 16109
rect 20290 15415 20414 15443
rect 20386 13667 20414 15415
rect 21250 14555 21278 16081
rect 21250 14527 21374 14555
rect 20962 13787 20990 14333
rect 20290 13639 20414 13667
rect 19522 12825 19646 12853
rect 19186 12159 19262 12187
rect 19042 11965 19070 12113
rect 18946 11937 19070 11965
rect 18274 11789 18398 11817
rect 18370 11225 18398 11789
rect 18274 11197 18398 11225
rect 18946 11225 18974 11937
rect 18946 11197 19166 11225
rect 18274 11049 18302 11197
rect 19138 10901 19166 11197
rect 17890 10827 18014 10855
rect 16450 10161 16574 10189
rect 16450 9597 16478 10161
rect 16450 9569 16574 9597
rect 16162 9495 16286 9523
rect 13378 8459 13502 8487
rect 13378 8237 13406 8459
rect 14914 8311 15134 8339
rect 11938 7571 12062 7599
rect 9922 6905 10046 6933
rect 9058 6017 9134 6045
rect 9106 5601 9134 6017
rect 9250 5647 9278 6239
rect 9106 5573 9182 5601
rect 8770 4121 8798 5083
rect 9154 4315 9182 5573
rect 9634 5009 9662 6831
rect 9634 4981 9758 5009
rect 9730 4713 9758 4981
rect 9634 4685 9758 4713
rect 7906 3723 8222 3751
rect 8674 4093 8798 4121
rect 6082 2539 6110 3011
rect 5602 2465 6014 2493
rect 4930 1827 4958 2123
rect 4930 1799 5054 1827
rect 34 985 158 1013
rect 34 51 62 985
rect 3586 911 3614 1207
rect 5026 1161 5054 1799
rect 5986 1577 6014 2465
rect 6178 1873 6206 2345
rect 6658 1873 6686 2937
rect 6850 2909 6878 3455
rect 7042 1725 7070 2123
rect 7906 1651 7934 3723
rect 8674 2937 8702 4093
rect 9634 4047 9662 4685
rect 9634 4019 9758 4047
rect 9730 3871 9758 4019
rect 8674 2909 8798 2937
rect 8674 2243 8702 2909
rect 9058 2567 9086 2937
rect 9922 2909 9950 6905
rect 10402 5129 10430 5675
rect 10594 4981 10622 6859
rect 10690 4491 10718 5453
rect 10690 4463 10814 4491
rect 8866 2539 9086 2567
rect 8866 1873 8894 2539
rect 9154 2391 9182 2789
rect 10306 1799 10334 4417
rect 10882 4343 10910 5527
rect 11074 5203 11102 6267
rect 11554 5647 11582 7007
rect 11938 5869 11966 7571
rect 12322 4537 12350 7673
rect 12994 6831 13022 7673
rect 13090 5869 13118 7007
rect 13282 6979 13310 7451
rect 13762 7201 13790 7673
rect 14050 6489 14078 7451
rect 13954 6461 14078 6489
rect 13954 5823 13982 6461
rect 13954 5795 14078 5823
rect 12706 5083 12734 5527
rect 12898 5203 12926 5675
rect 12706 5055 12830 5083
rect 10690 4315 10910 4343
rect 12706 4343 12734 5055
rect 12706 4315 12926 4343
rect 10690 3159 10718 4315
rect 10978 3205 11006 4269
rect 10690 3131 10910 3159
rect 4930 1133 5054 1161
rect 4930 985 4958 1133
rect 10690 1059 10718 2937
rect 10882 2539 10910 3131
rect 12706 2539 12734 4315
rect 13090 3205 13118 4491
rect 13186 1059 13214 1753
rect 13474 1207 13502 5009
rect 13858 2983 13886 5675
rect 14050 5203 14078 5795
rect 14242 4241 14270 7599
rect 14338 7201 14366 8191
rect 14530 6535 14558 7451
rect 14722 7155 14750 8117
rect 14914 7571 14942 8311
rect 15010 7867 15038 8265
rect 15106 8237 15134 8311
rect 15202 7793 15230 9005
rect 15586 8977 15614 9449
rect 16258 9153 16286 9495
rect 16066 9125 16286 9153
rect 16066 8413 16094 9125
rect 16546 8857 16574 9569
rect 16354 8829 16574 8857
rect 16066 8385 16286 8413
rect 15394 7747 15422 8265
rect 16258 8237 16286 8385
rect 15394 7719 15518 7747
rect 15202 7201 15230 7451
rect 15490 7155 15518 7719
rect 14722 7127 14846 7155
rect 14530 3825 14558 6415
rect 14818 6193 14846 7127
rect 15394 7127 15518 7155
rect 15394 6535 15422 7127
rect 14722 6165 14846 6193
rect 14722 5869 14750 6165
rect 15874 5675 15902 6933
rect 15490 5647 15902 5675
rect 16354 5647 16382 8829
rect 16450 8237 16478 8783
rect 16834 8533 16862 9449
rect 17314 9051 17342 9597
rect 17506 8533 17534 10115
rect 17602 8117 17630 8265
rect 17506 8089 17630 8117
rect 16642 5675 16670 7747
rect 17506 7599 17534 8089
rect 17506 7571 17630 7599
rect 17602 7423 17630 7571
rect 17794 7201 17822 10337
rect 17986 9051 18014 10827
rect 18946 10309 18974 10781
rect 19234 10309 19262 12159
rect 18178 9865 18206 10115
rect 19330 9865 19358 10411
rect 19522 9791 19550 12825
rect 19906 10753 19934 12113
rect 20290 11521 20318 13639
rect 21250 13149 21278 14407
rect 21346 14305 21374 14527
rect 21154 13121 21278 13149
rect 21154 12557 21182 13121
rect 21154 12529 21278 12557
rect 21346 12529 21374 13075
rect 21538 12973 21566 16969
rect 21634 16183 21662 16775
rect 21922 16377 21950 17635
rect 23074 16997 23102 17663
rect 23074 16969 23198 16997
rect 22978 16775 23006 16923
rect 22882 16747 23006 16775
rect 22882 16257 22910 16747
rect 22882 16229 23006 16257
rect 21634 16155 21758 16183
rect 21730 14555 21758 16155
rect 22978 16081 23006 16229
rect 23170 16183 23198 16969
rect 23746 16525 23774 17589
rect 24034 16895 24062 20919
rect 24130 20891 24350 20919
rect 24226 19041 24254 19439
rect 24322 19189 24350 20891
rect 24322 17857 24350 18255
rect 24226 17191 24254 17589
rect 24706 16553 24734 32315
rect 25186 23111 25214 26321
rect 25474 25035 25502 28319
rect 26050 25063 26078 27653
rect 26530 25701 26558 28393
rect 26434 25183 26462 25581
rect 26050 25035 26366 25063
rect 25858 24517 25886 24767
rect 25378 21631 25406 23139
rect 25858 22519 25886 22769
rect 26050 22325 26078 25035
rect 25762 22297 26078 22325
rect 25474 18301 25502 21659
rect 25762 21511 25790 22297
rect 25762 21483 25886 21511
rect 25858 21039 25886 21483
rect 26050 20817 26078 22251
rect 26338 22223 26366 24397
rect 26530 22741 26558 24989
rect 26722 24175 26750 24323
rect 26722 24147 26846 24175
rect 26818 23509 26846 24147
rect 26722 23481 26846 23509
rect 26722 21733 26750 23481
rect 27106 22991 27134 23139
rect 27010 22963 27134 22991
rect 27010 22177 27038 22963
rect 27298 22547 27326 25433
rect 27682 25211 27710 28097
rect 28450 27847 28478 28393
rect 29122 26515 29150 27727
rect 29890 27283 29918 27431
rect 29794 27255 29918 27283
rect 27682 25183 27806 25211
rect 28546 24841 28574 26395
rect 28450 24813 28574 24841
rect 28450 23139 28478 24813
rect 28450 23111 28574 23139
rect 27490 22843 27518 22991
rect 27490 22815 27614 22843
rect 27298 22519 27422 22547
rect 27010 22149 27134 22177
rect 26722 21705 26846 21733
rect 25858 19707 25886 20771
rect 26050 18329 26078 18477
rect 25954 18301 26078 18329
rect 24898 17857 24926 18255
rect 25954 17737 25982 18301
rect 25954 17709 26078 17737
rect 25474 17191 25502 17441
rect 24706 16525 24830 16553
rect 23074 16155 23198 16183
rect 23074 16035 23102 16155
rect 22978 16007 23102 16035
rect 21634 14527 21758 14555
rect 21922 14527 21950 15665
rect 22978 14971 23006 16007
rect 23842 15119 23870 16331
rect 25858 15193 25886 16109
rect 26050 15813 26078 17709
rect 26242 17561 26270 21585
rect 26530 17783 26558 21659
rect 26818 21141 26846 21705
rect 26722 21113 26846 21141
rect 26722 20965 26750 21113
rect 26050 15785 26270 15813
rect 26338 15563 26366 16331
rect 26626 16109 26654 18107
rect 26434 16081 26654 16109
rect 21634 14407 21662 14527
rect 21634 14379 21854 14407
rect 21730 13417 21758 14111
rect 21826 13861 21854 14379
rect 20674 11715 20702 12335
rect 21058 11863 21086 12335
rect 21250 11715 21278 12529
rect 22306 12409 22334 14777
rect 24610 14527 24638 14925
rect 25378 14527 25406 14925
rect 22978 13001 23006 14333
rect 23746 13713 23774 14407
rect 22978 12973 23198 13001
rect 22978 12529 23006 12927
rect 23170 12483 23198 12973
rect 24226 12631 24254 12779
rect 23074 12455 23198 12483
rect 24034 12603 24254 12631
rect 22306 12381 22430 12409
rect 20194 11493 20318 11521
rect 18274 9199 18302 9671
rect 18082 7081 18110 8783
rect 18466 8459 18494 9005
rect 18946 8311 18974 9523
rect 18274 7821 18302 8265
rect 18274 7793 18398 7821
rect 17986 7053 18110 7081
rect 17698 6535 17726 7007
rect 16642 5647 16766 5675
rect 15106 4315 15134 5453
rect 14530 3797 14654 3825
rect 14338 3529 14366 3677
rect 14242 3501 14366 3529
rect 14242 2493 14270 3501
rect 14242 2465 14366 2493
rect 14338 2317 14366 2465
rect 14530 2391 14558 3797
rect 14818 3723 14846 4121
rect 14722 2391 14750 2789
rect 15490 2493 15518 5647
rect 15778 2539 15806 5601
rect 16258 5055 16286 5453
rect 16738 5203 16766 5647
rect 17314 4907 17342 5675
rect 17698 4981 17726 5453
rect 17986 4935 18014 7053
rect 18370 7007 18398 7793
rect 19234 7525 19262 9671
rect 19522 8533 19550 9671
rect 20194 9597 20222 11493
rect 20386 11197 20414 11447
rect 21730 11299 21758 11447
rect 21634 11271 21758 11299
rect 20482 9643 20510 10781
rect 20194 9569 20318 9597
rect 20098 9199 20126 9449
rect 20290 9421 20318 9569
rect 19234 7497 19358 7525
rect 18274 6979 18398 7007
rect 17986 4907 18110 4935
rect 18082 4463 18110 4907
rect 18274 4537 18302 6979
rect 19138 6933 19166 7451
rect 19042 6905 19166 6933
rect 19042 6415 19070 6905
rect 19330 6859 19358 7497
rect 19522 6979 19550 8339
rect 19282 6831 19358 6859
rect 19042 6387 19166 6415
rect 19042 5647 19070 6267
rect 19138 6165 19166 6387
rect 19282 6119 19310 6831
rect 19714 6387 19742 6785
rect 19234 6091 19310 6119
rect 19234 5055 19262 6091
rect 19234 4787 19262 4935
rect 19138 4759 19262 4787
rect 15490 2465 15614 2493
rect 14626 985 14654 1679
rect 15586 1207 15614 2465
rect 16450 1133 16478 4269
rect 16834 3871 16862 4269
rect 17890 3057 17918 3455
rect 18082 2909 18110 3825
rect 18274 3649 18302 4121
rect 18658 3205 18686 4343
rect 19138 4269 19166 4759
rect 18850 3649 18878 4269
rect 19138 4241 19262 4269
rect 19234 4093 19262 4241
rect 19426 3797 19454 6341
rect 19714 5203 19742 5601
rect 20098 4981 20126 8487
rect 20482 7821 20510 9153
rect 20674 8533 20702 9597
rect 20386 7793 20510 7821
rect 21058 7793 21086 10929
rect 21634 10411 21662 11271
rect 21634 10383 21758 10411
rect 21730 10235 21758 10383
rect 21442 8311 21470 9227
rect 20386 4537 20414 7793
rect 19810 3871 19838 4269
rect 19426 2345 19454 3677
rect 19426 2317 19550 2345
rect 20386 2317 20414 3751
rect 18178 1207 18206 2271
rect 20098 1873 20126 2271
rect 20674 1207 20702 7747
rect 21634 7645 21662 8783
rect 21730 8533 21758 9005
rect 21922 8533 21950 11817
rect 22306 11225 22334 12335
rect 22402 11641 22430 12381
rect 22306 11197 22430 11225
rect 22210 8783 22238 9597
rect 22306 9569 22334 10115
rect 22498 9717 22526 11743
rect 23074 10383 23102 12455
rect 23554 11863 23582 12113
rect 23266 11197 23294 11447
rect 23266 9643 23294 10115
rect 23074 8903 23102 9449
rect 23458 9375 23486 10411
rect 23746 10161 23774 12113
rect 24034 11373 24062 12603
rect 24034 11345 24254 11373
rect 24034 10309 24062 11225
rect 23650 9569 23678 10115
rect 23842 9865 23870 10263
rect 23458 9347 23678 9375
rect 23650 8977 23678 9347
rect 24226 9079 24254 11345
rect 24322 10975 24350 14111
rect 24994 11197 25022 12409
rect 25474 12233 25502 14333
rect 26434 13741 26462 14999
rect 26722 13861 26750 16109
rect 27106 14925 27134 22149
rect 27298 21853 27326 22251
rect 27586 21807 27614 22815
rect 27490 21779 27614 21807
rect 27490 20993 27518 21779
rect 27874 21557 27902 22991
rect 28354 22371 28382 22991
rect 28546 22297 28574 23111
rect 27394 20965 27518 20993
rect 27394 19809 27422 20965
rect 27682 19855 27710 20919
rect 27394 19781 27806 19809
rect 27298 17709 27326 18107
rect 27010 14897 27134 14925
rect 27010 14185 27038 14897
rect 27010 14157 27134 14185
rect 26434 13713 26558 13741
rect 25666 12307 25694 12779
rect 25858 12529 25886 13593
rect 26050 11817 26078 13667
rect 25954 11789 26078 11817
rect 25954 11077 25982 11789
rect 25954 11049 26078 11077
rect 26050 10531 26078 11049
rect 25090 9199 25118 9449
rect 25378 9199 25406 9597
rect 26242 9125 26270 13445
rect 26434 12899 26462 13713
rect 26626 12973 26654 13445
rect 26434 10457 26462 10781
rect 24130 9051 24254 9079
rect 22210 8755 22334 8783
rect 22306 8533 22334 8755
rect 21826 6535 21854 7673
rect 22114 7451 22142 8117
rect 22978 7747 23006 8339
rect 22978 7719 23102 7747
rect 22114 7423 22334 7451
rect 22306 6535 22334 7423
rect 22786 7201 22814 7673
rect 23074 7155 23102 7719
rect 22978 7127 23102 7155
rect 21058 5203 21086 6341
rect 22306 5721 22334 6119
rect 22786 5203 22814 5601
rect 21058 3899 21086 4121
rect 20962 3871 21086 3899
rect 20962 2789 20990 3871
rect 20962 2761 21086 2789
rect 21058 1235 21086 2761
rect 21154 2539 21182 5009
rect 21442 2983 21470 5009
rect 22690 3131 22718 3455
rect 22786 3205 22814 3603
rect 22978 3205 23006 7127
rect 23458 6979 23486 8413
rect 23554 8311 23582 8783
rect 23074 6415 23102 6933
rect 24226 6859 24254 8931
rect 24706 8533 24734 8783
rect 25474 8311 25502 8931
rect 25666 8533 25694 9079
rect 25474 7053 25502 8117
rect 24130 6831 24254 6859
rect 23074 6387 23486 6415
rect 23458 4537 23486 6387
rect 23650 4491 23678 5157
rect 23746 4981 23774 6119
rect 24130 5823 24158 6831
rect 25186 6785 25214 6933
rect 24418 6119 24446 6785
rect 24322 6091 24446 6119
rect 25090 6757 25214 6785
rect 24322 5869 24350 6091
rect 25090 5823 25118 6757
rect 24130 5795 24254 5823
rect 25090 5795 25214 5823
rect 24226 5203 24254 5795
rect 25186 5647 25214 5795
rect 25378 5721 25406 7007
rect 26242 6267 26270 6415
rect 26146 6239 26270 6267
rect 26146 5527 26174 6239
rect 26434 5573 26462 8931
rect 26722 7201 26750 8783
rect 26146 5499 26270 5527
rect 26242 5203 26270 5499
rect 26626 5453 26654 6119
rect 26530 5425 26654 5453
rect 26530 4935 26558 5425
rect 26722 4981 26750 5453
rect 26530 4907 26654 4935
rect 23458 4463 23678 4491
rect 23170 3205 23198 3677
rect 23458 2493 23486 4463
rect 26626 4389 26654 4907
rect 23650 4121 23678 4269
rect 23650 4093 23774 4121
rect 23746 3159 23774 4093
rect 24514 3455 24542 4269
rect 25954 3649 25982 4121
rect 26146 3797 26174 4269
rect 24514 3427 24734 3455
rect 24706 3205 24734 3427
rect 23362 2465 23486 2493
rect 23650 3131 23774 3159
rect 23362 1901 23390 2465
rect 23650 2123 23678 3131
rect 26818 2317 26846 2937
rect 27010 2243 27038 3011
rect 27106 2539 27134 14157
rect 27298 14037 27326 14851
rect 27394 14083 27422 14777
rect 27586 14555 27614 18329
rect 27778 17783 27806 19781
rect 28162 18995 28190 19069
rect 28162 18967 28286 18995
rect 28258 18477 28286 18967
rect 28450 18847 28478 20993
rect 28738 18921 28766 24767
rect 29026 24443 29054 26247
rect 29794 24027 29822 27255
rect 29794 23999 29918 24027
rect 29890 23851 29918 23999
rect 30082 23731 30110 31205
rect 32002 31177 32030 32583
rect 31522 31103 32064 31131
rect 30946 27579 30974 29651
rect 30946 27551 31070 27579
rect 31042 26839 31070 27551
rect 30946 26811 31070 26839
rect 30946 25063 30974 26811
rect 30946 25035 31070 25063
rect 30562 24471 30590 24989
rect 29986 23703 30110 23731
rect 30274 24443 30590 24471
rect 29026 21039 29054 23583
rect 29122 21807 29150 22103
rect 29122 21779 29342 21807
rect 28930 19041 28958 20919
rect 29314 20845 29342 21779
rect 29122 20817 29342 20845
rect 29122 20475 29150 20817
rect 29122 20447 29246 20475
rect 29218 19513 29246 20447
rect 29122 19485 29246 19513
rect 28738 18893 28862 18921
rect 28450 18819 28574 18847
rect 28162 18449 28286 18477
rect 27586 14527 27710 14555
rect 27682 14305 27710 14527
rect 27874 14231 27902 17737
rect 28162 17515 28190 18449
rect 28450 18375 28478 18773
rect 28546 18329 28574 18819
rect 28450 18301 28574 18329
rect 28162 17487 28286 17515
rect 28258 16969 28286 17487
rect 28450 17043 28478 18301
rect 28834 18255 28862 18893
rect 28738 18227 28862 18255
rect 28258 15711 28286 16775
rect 28450 14379 28478 15443
rect 27298 14009 27422 14037
rect 27394 13593 27422 14009
rect 27394 13565 27518 13593
rect 27394 9643 27422 13565
rect 27682 9865 27710 10263
rect 27874 9791 27902 12927
rect 28066 12529 28094 13001
rect 28258 12973 28286 13593
rect 27778 8829 27806 9597
rect 28258 8977 28286 12335
rect 28546 11715 28574 12779
rect 28738 9745 28766 18227
rect 29122 12483 29150 19485
rect 29410 18107 29438 19069
rect 29410 18079 29534 18107
rect 29506 17857 29534 18079
rect 29410 15711 29438 16257
rect 29122 12455 29246 12483
rect 28930 11863 28958 12409
rect 29218 11817 29246 12455
rect 28642 9717 28766 9745
rect 29122 11789 29246 11817
rect 29122 9745 29150 11789
rect 29602 10559 29630 21437
rect 29986 20401 30014 23703
rect 30274 23555 30302 24443
rect 30754 24397 30782 24915
rect 30658 24369 30782 24397
rect 30658 23879 30686 24369
rect 31042 24249 31070 25035
rect 30466 23851 30686 23879
rect 30946 24221 31070 24249
rect 29890 20373 30014 20401
rect 29890 17071 29918 20373
rect 30274 20327 30302 23435
rect 30466 23361 30494 23851
rect 30466 23333 30686 23361
rect 30658 20845 30686 23333
rect 30946 21659 30974 24221
rect 31234 21705 31262 26765
rect 30946 21631 31070 21659
rect 30178 20299 30302 20327
rect 30562 20817 30686 20845
rect 30178 17145 30206 20299
rect 30562 20179 30590 20817
rect 30562 20151 30686 20179
rect 30658 19633 30686 20151
rect 30754 19291 30782 20845
rect 31042 19707 31070 21631
rect 31138 20697 31166 20845
rect 31138 20669 31262 20697
rect 31234 19587 31262 20669
rect 30658 19263 30782 19291
rect 30178 17117 30398 17145
rect 29890 17043 30110 17071
rect 29890 14527 29918 16923
rect 30082 15637 30110 17043
rect 30370 16183 30398 17117
rect 30274 16155 30398 16183
rect 29602 10531 29822 10559
rect 29122 9717 29246 9745
rect 28642 8931 28670 9717
rect 28930 8977 28958 9671
rect 29218 8931 29246 9717
rect 29506 9643 29534 10485
rect 29794 9597 29822 10531
rect 28642 8903 28766 8931
rect 27682 4861 27710 7007
rect 28738 5869 28766 8903
rect 29122 8903 29246 8931
rect 29602 9569 29822 9597
rect 29122 6091 29150 8903
rect 29602 8533 29630 9569
rect 27586 4833 27710 4861
rect 27586 3159 27614 4833
rect 27586 3131 27710 3159
rect 27682 2983 27710 3131
rect 27874 2909 27902 5083
rect 28258 3057 28286 4121
rect 29602 3205 29630 4343
rect 30274 2909 30302 16155
rect 30658 15637 30686 19263
rect 30946 17191 30974 19587
rect 31138 19559 31262 19587
rect 30850 16229 30878 16775
rect 30946 15295 30974 15443
rect 30850 15267 30974 15295
rect 30850 13001 30878 15267
rect 30850 12973 30974 13001
rect 30946 12825 30974 12973
rect 31138 12705 31166 19559
rect 31330 18329 31358 19439
rect 31522 19143 31550 31103
rect 31906 29623 32064 29651
rect 31967 28143 32064 28171
rect 32002 26737 32030 28143
rect 31906 26663 32064 26691
rect 31906 26367 31934 26663
rect 31810 25183 32064 25211
rect 31810 25109 31838 25183
rect 31906 23703 32064 23731
rect 31618 22815 31742 22843
rect 31714 22251 31742 22815
rect 31714 22223 32064 22251
rect 31906 20743 32064 20771
rect 31967 19263 32064 19291
rect 31522 19115 31646 19143
rect 31618 18551 31646 19115
rect 32002 18819 32030 19263
rect 31522 18523 31646 18551
rect 31522 18375 31550 18523
rect 31330 18301 31454 18329
rect 31042 12677 31166 12705
rect 31042 10411 31070 12677
rect 31330 10457 31358 18107
rect 31426 17737 31454 18301
rect 31906 17783 32064 17811
rect 31426 17709 31646 17737
rect 31618 16849 31646 17709
rect 31522 16821 31646 16849
rect 31522 16479 31550 16821
rect 31522 16451 31646 16479
rect 31618 15517 31646 16451
rect 32002 16331 32030 17589
rect 31967 16303 32064 16331
rect 31522 15489 31646 15517
rect 31522 15147 31550 15489
rect 31522 15119 31646 15147
rect 31618 14185 31646 15119
rect 32002 14851 32030 15221
rect 31967 14823 32064 14851
rect 31522 14157 31646 14185
rect 31522 13815 31550 14157
rect 31522 13787 31646 13815
rect 31618 12853 31646 13787
rect 32002 13371 32030 13889
rect 31967 13343 32064 13371
rect 31522 12825 31646 12853
rect 31522 12483 31550 12825
rect 31522 12455 31646 12483
rect 31618 11521 31646 12455
rect 32002 11891 32030 12853
rect 31967 11863 32064 11891
rect 31522 11493 31646 11521
rect 31522 11151 31550 11493
rect 31522 11123 31646 11151
rect 31618 10411 31646 11123
rect 32002 10411 32030 10485
rect 31042 10383 31166 10411
rect 31618 10383 31934 10411
rect 31967 10383 32064 10411
rect 23650 2095 23774 2123
rect 23362 1873 23486 1901
rect 20962 1207 21086 1235
rect 20962 985 20990 1207
rect 21250 985 21278 1605
rect 23458 1059 23486 1873
rect 23650 1059 23678 2095
rect 27106 1873 27134 2271
rect 24130 985 24158 1679
rect 31138 51 31166 10383
rect 31906 8931 31934 10383
rect 31906 8903 32064 8931
rect 31810 7451 31838 8561
rect 31810 7423 32064 7451
rect 31906 5971 31934 6119
rect 31906 5943 32064 5971
rect 32002 4491 32030 5897
rect 31967 4463 32064 4491
rect 31906 2983 32064 3011
rect 31906 2909 31934 2983
rect 32002 1531 32030 2567
rect 31967 1503 32064 1531
rect 0 23 97 51
rect 31138 23 32064 51
<< metal3 >>
rect 400 0 600 32634
rect 1600 0 1800 32634
rect 2800 0 3000 32634
rect 4000 0 4200 32634
rect 5200 0 5400 32634
rect 6400 0 6600 32634
rect 7600 0 7800 32634
rect 8800 0 9000 32634
rect 10000 0 10200 32634
rect 11200 0 11400 32634
rect 12400 0 12600 32634
rect 13600 0 13800 32634
rect 14800 0 15000 32634
rect 16000 0 16200 32634
rect 17200 0 17400 32634
rect 18400 0 18600 32634
rect 19600 0 19800 32634
rect 20800 0 21000 32634
rect 22000 0 22200 32634
rect 23200 0 23400 32634
rect 24400 0 24600 32634
rect 25600 0 25800 32634
rect 26800 0 27000 32634
rect 28000 0 28200 32634
rect 29200 0 29400 32634
rect 30400 0 30600 32634
rect 31600 0 31800 32634
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_356
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_713
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_345
timestamp 1626908933
transform 1 0 0 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_356
timestamp 1626908933
transform 1 0 0 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_946
timestamp 1626908933
transform 1 0 0 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_957
timestamp 1626908933
transform 1 0 0 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_648
timestamp 1626908933
transform 1 0 192 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1639
timestamp 1626908933
transform 1 0 192 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_335
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_983
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_335
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_983
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_699
timestamp 1626908933
transform 1 0 768 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_721
timestamp 1626908933
transform 1 0 192 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1421
timestamp 1626908933
transform 1 0 768 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1443
timestamp 1626908933
transform 1 0 192 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_595
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1193
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_628
timestamp 1626908933
transform 1 0 960 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1619
timestamp 1626908933
transform 1 0 960 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_355
timestamp 1626908933
transform 1 0 1536 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_956
timestamp 1626908933
transform 1 0 1536 0 1 0
box -38 -49 230 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_26
timestamp 1626908933
transform 1 0 1700 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_53
timestamp 1626908933
transform 1 0 1700 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_26
timestamp 1626908933
transform 1 0 1700 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_53
timestamp 1626908933
transform 1 0 1700 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_688
timestamp 1626908933
transform 1 0 1440 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1410
timestamp 1626908933
transform 1 0 1440 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_584
timestamp 1626908933
transform 1 0 1056 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1182
timestamp 1626908933
transform 1 0 1056 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_342
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_355
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_699
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_712
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_358
timestamp 1626908933
transform 1 0 2304 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_959
timestamp 1626908933
transform 1 0 2304 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_627
timestamp 1626908933
transform 1 0 2208 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1618
timestamp 1626908933
transform 1 0 2208 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_665
timestamp 1626908933
transform 1 0 1728 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1387
timestamp 1626908933
transform 1 0 1728 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1638
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_647
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1146
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_548
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1380
timestamp 1626908933
transform 1 0 2688 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_658
timestamp 1626908933
transform 1 0 2688 0 1 0
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_959
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_311
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_959
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_311
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_12
timestamp 1626908933
transform 1 0 2976 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_4
timestamp 1626908933
transform 1 0 2976 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1139
timestamp 1626908933
transform 1 0 3456 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_541
timestamp 1626908933
transform 1 0 3456 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_344
timestamp 1626908933
transform 1 0 3648 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_354
timestamp 1626908933
transform 1 0 3840 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_945
timestamp 1626908933
transform 1 0 3648 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_955
timestamp 1626908933
transform 1 0 3840 0 1 0
box -38 -49 230 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_25
timestamp 1626908933
transform 1 0 4100 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_52
timestamp 1626908933
transform 1 0 4100 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_25
timestamp 1626908933
transform 1 0 4100 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_52
timestamp 1626908933
transform 1 0 4100 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_635
timestamp 1626908933
transform 1 0 4032 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1357
timestamp 1626908933
transform 1 0 4032 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_529
timestamp 1626908933
transform 1 0 3840 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1127
timestamp 1626908933
transform 1 0 3840 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_6
timestamp 1626908933
transform 1 0 4224 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_14
timestamp 1626908933
transform 1 0 4224 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_646
timestamp 1626908933
transform 1 0 4800 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1637
timestamp 1626908933
transform 1 0 4800 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1640
timestamp 1626908933
transform 1 0 4896 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_649
timestamp 1626908933
transform 1 0 4896 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_711
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_354
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_935
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_287
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_935
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_287
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_954
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_353
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_612
timestamp 1626908933
transform 1 0 5280 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_613
timestamp 1626908933
transform 1 0 5280 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1334
timestamp 1626908933
transform 1 0 5280 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1335
timestamp 1626908933
transform 1 0 5280 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_512
timestamp 1626908933
transform 1 0 4896 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1110
timestamp 1626908933
transform 1 0 4896 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1094
timestamp 1626908933
transform 1 0 6048 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1093
timestamp 1626908933
transform 1 0 6048 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_496
timestamp 1626908933
transform 1 0 6048 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_495
timestamp 1626908933
transform 1 0 6048 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_626
timestamp 1626908933
transform 1 0 6432 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_645
timestamp 1626908933
transform 1 0 6432 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1617
timestamp 1626908933
transform 1 0 6432 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1636
timestamp 1626908933
transform 1 0 6432 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_24
timestamp 1626908933
transform 1 0 6500 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_51
timestamp 1626908933
transform 1 0 6500 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_24
timestamp 1626908933
transform 1 0 6500 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_51
timestamp 1626908933
transform 1 0 6500 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_584
timestamp 1626908933
transform 1 0 6528 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_585
timestamp 1626908933
transform 1 0 6528 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1306
timestamp 1626908933
transform 1 0 6528 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1307
timestamp 1626908933
transform 1 0 6528 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1648
timestamp 1626908933
transform 1 0 7392 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1641
timestamp 1626908933
transform 1 0 7392 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1635
timestamp 1626908933
transform 1 0 7296 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1616
timestamp 1626908933
transform 1 0 7296 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_657
timestamp 1626908933
transform 1 0 7392 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_650
timestamp 1626908933
transform 1 0 7392 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_644
timestamp 1626908933
transform 1 0 7296 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_625
timestamp 1626908933
transform 1 0 7296 0 -1 1332
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_911
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_263
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_911
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_263
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_710
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_698
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_353
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_341
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_953
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_944
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_352
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_343
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_624
timestamp 1626908933
transform 1 0 7776 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_643
timestamp 1626908933
transform 1 0 7776 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1615
timestamp 1626908933
transform 1 0 7776 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1634
timestamp 1626908933
transform 1 0 7776 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_562
timestamp 1626908933
transform 1 0 7872 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_563
timestamp 1626908933
transform 1 0 7872 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1284
timestamp 1626908933
transform 1 0 7872 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1285
timestamp 1626908933
transform 1 0 7872 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_623
timestamp 1626908933
transform 1 0 8640 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_642
timestamp 1626908933
transform 1 0 8640 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1614
timestamp 1626908933
transform 1 0 8640 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1633
timestamp 1626908933
transform 1 0 8640 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_23
timestamp 1626908933
transform 1 0 8900 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_50
timestamp 1626908933
transform 1 0 8900 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_23
timestamp 1626908933
transform 1 0 8900 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_50
timestamp 1626908933
transform 1 0 8900 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_542
timestamp 1626908933
transform 1 0 9120 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_543
timestamp 1626908933
transform 1 0 9120 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1264
timestamp 1626908933
transform 1 0 9120 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1265
timestamp 1626908933
transform 1 0 9120 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_451
timestamp 1626908933
transform 1 0 8736 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_452
timestamp 1626908933
transform 1 0 8736 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1049
timestamp 1626908933
transform 1 0 8736 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1050
timestamp 1626908933
transform 1 0 8736 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1642
timestamp 1626908933
transform 1 0 9888 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_651
timestamp 1626908933
transform 1 0 9888 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_943
timestamp 1626908933
transform 1 0 9888 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_342
timestamp 1626908933
transform 1 0 9888 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_709
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_352
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_239
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_887
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_239
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_887
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_522
timestamp 1626908933
transform 1 0 10464 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_523
timestamp 1626908933
transform 1 0 10464 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1244
timestamp 1626908933
transform 1 0 10464 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1245
timestamp 1626908933
transform 1 0 10464 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_428
timestamp 1626908933
transform 1 0 10080 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_429
timestamp 1626908933
transform 1 0 10080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1026
timestamp 1626908933
transform 1 0 10080 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1027
timestamp 1626908933
transform 1 0 10080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_622
timestamp 1626908933
transform 1 0 11232 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_641
timestamp 1626908933
transform 1 0 11232 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1613
timestamp 1626908933
transform 1 0 11232 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1632
timestamp 1626908933
transform 1 0 11232 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_22
timestamp 1626908933
transform 1 0 11300 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_49
timestamp 1626908933
transform 1 0 11300 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_22
timestamp 1626908933
transform 1 0 11300 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_49
timestamp 1626908933
transform 1 0 11300 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_489
timestamp 1626908933
transform 1 0 11712 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_490
timestamp 1626908933
transform 1 0 11712 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1211
timestamp 1626908933
transform 1 0 11712 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1212
timestamp 1626908933
transform 1 0 11712 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_402
timestamp 1626908933
transform 1 0 11328 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_403
timestamp 1626908933
transform 1 0 11328 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1000
timestamp 1626908933
transform 1 0 11328 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1001
timestamp 1626908933
transform 1 0 11328 0 1 0
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_863
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_215
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_863
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_215
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_708
timestamp 1626908933
transform 1 0 12480 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_697
timestamp 1626908933
transform 1 0 12480 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_351
timestamp 1626908933
transform 1 0 12480 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_340
timestamp 1626908933
transform 1 0 12480 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_942
timestamp 1626908933
transform 1 0 12576 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_341
timestamp 1626908933
transform 1 0 12576 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_368
timestamp 1626908933
transform 1 0 12576 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_966
timestamp 1626908933
transform 1 0 12576 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_941
timestamp 1626908933
transform 1 0 13440 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_340
timestamp 1626908933
transform 1 0 13440 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_965
timestamp 1626908933
transform 1 0 12768 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_367
timestamp 1626908933
transform 1 0 12768 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1189
timestamp 1626908933
transform 1 0 12960 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_467
timestamp 1626908933
transform 1 0 12960 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_81
timestamp 1626908933
transform 1 0 13152 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_20
timestamp 1626908933
transform 1 0 13152 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_640
timestamp 1626908933
transform 1 0 13728 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1631
timestamp 1626908933
transform 1 0 13728 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_21
timestamp 1626908933
transform 1 0 13700 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_48
timestamp 1626908933
transform 1 0 13700 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_21
timestamp 1626908933
transform 1 0 13700 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_48
timestamp 1626908933
transform 1 0 13700 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_450
timestamp 1626908933
transform 1 0 13632 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1172
timestamp 1626908933
transform 1 0 13632 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_347
timestamp 1626908933
transform 1 0 13824 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_945
timestamp 1626908933
transform 1 0 13824 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1612
timestamp 1626908933
transform 1 0 14400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_621
timestamp 1626908933
transform 1 0 14400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_936
timestamp 1626908933
transform 1 0 14496 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_338
timestamp 1626908933
transform 1 0 14496 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1157
timestamp 1626908933
transform 1 0 14208 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_435
timestamp 1626908933
transform 1 0 14208 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_350
timestamp 1626908933
transform 1 0 14976 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_707
timestamp 1626908933
transform 1 0 14976 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_191
timestamp 1626908933
transform 1 0 14900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_839
timestamp 1626908933
transform 1 0 14900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_191
timestamp 1626908933
transform 1 0 14900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_839
timestamp 1626908933
transform 1 0 14900 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_639
timestamp 1626908933
transform 1 0 15456 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1630
timestamp 1626908933
transform 1 0 15456 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_423
timestamp 1626908933
transform 1 0 14880 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1145
timestamp 1626908933
transform 1 0 14880 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_326
timestamp 1626908933
transform 1 0 15072 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_924
timestamp 1626908933
transform 1 0 15072 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_620
timestamp 1626908933
transform 1 0 15648 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1611
timestamp 1626908933
transform 1 0 15648 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_24
timestamp 1626908933
transform -1 0 16032 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_86
timestamp 1626908933
transform -1 0 16032 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_339
timestamp 1626908933
transform 1 0 16032 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_940
timestamp 1626908933
transform 1 0 16032 0 -1 1332
box -38 -49 230 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_20
timestamp 1626908933
transform 1 0 16100 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_47
timestamp 1626908933
transform 1 0 16100 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_20
timestamp 1626908933
transform 1 0 16100 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_47
timestamp 1626908933
transform 1 0 16100 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_396
timestamp 1626908933
transform 1 0 16224 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_418
timestamp 1626908933
transform 1 0 15552 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1118
timestamp 1626908933
transform 1 0 16224 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1140
timestamp 1626908933
transform 1 0 15552 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_299
timestamp 1626908933
transform 1 0 16320 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_897
timestamp 1626908933
transform 1 0 16320 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_619
timestamp 1626908933
transform 1 0 16992 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1610
timestamp 1626908933
transform 1 0 16992 0 -1 1332
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_167
timestamp 1626908933
transform 1 0 17300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_815
timestamp 1626908933
transform 1 0 17300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_167
timestamp 1626908933
transform 1 0 17300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_815
timestamp 1626908933
transform 1 0 17300 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_388
timestamp 1626908933
transform 1 0 16704 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1110
timestamp 1626908933
transform 1 0 16704 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_284
timestamp 1626908933
transform 1 0 17088 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_882
timestamp 1626908933
transform 1 0 17088 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_339
timestamp 1626908933
transform 1 0 17472 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_349
timestamp 1626908933
transform 1 0 17472 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_696
timestamp 1626908933
transform 1 0 17472 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_706
timestamp 1626908933
transform 1 0 17472 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_638
timestamp 1626908933
transform 1 0 17568 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1629
timestamp 1626908933
transform 1 0 17568 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_637
timestamp 1626908933
transform 1 0 18048 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1628
timestamp 1626908933
transform 1 0 18048 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_365
timestamp 1626908933
transform 1 0 18144 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1087
timestamp 1626908933
transform 1 0 18144 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_277
timestamp 1626908933
transform 1 0 17664 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_875
timestamp 1626908933
transform 1 0 17664 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_9
timestamp 1626908933
transform 1 0 17568 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_61
timestamp 1626908933
transform 1 0 17568 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_16
timestamp 1626908933
transform 1 0 17952 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_78
timestamp 1626908933
transform 1 0 17952 0 -1 1332
box -38 -49 422 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_19
timestamp 1626908933
transform 1 0 18500 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_46
timestamp 1626908933
transform 1 0 18500 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_19
timestamp 1626908933
transform 1 0 18500 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_46
timestamp 1626908933
transform 1 0 18500 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_351
timestamp 1626908933
transform 1 0 18912 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_952
timestamp 1626908933
transform 1 0 18912 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_636
timestamp 1626908933
transform 1 0 19104 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1627
timestamp 1626908933
transform 1 0 19104 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_341
timestamp 1626908933
transform 1 0 18720 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1063
timestamp 1626908933
transform 1 0 18720 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_249
timestamp 1626908933
transform 1 0 18336 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_847
timestamp 1626908933
transform 1 0 18336 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1056
timestamp 1626908933
transform 1 0 19200 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_334
timestamp 1626908933
transform 1 0 19200 0 1 0
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_143
timestamp 1626908933
transform 1 0 19700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_791
timestamp 1626908933
transform 1 0 19700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_143
timestamp 1626908933
transform 1 0 19700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_791
timestamp 1626908933
transform 1 0 19700 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_348
timestamp 1626908933
transform 1 0 19968 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_705
timestamp 1626908933
transform 1 0 19968 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_338
timestamp 1626908933
transform 1 0 19872 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_939
timestamp 1626908933
transform 1 0 19872 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_313
timestamp 1626908933
transform 1 0 20064 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_314
timestamp 1626908933
transform 1 0 20064 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1035
timestamp 1626908933
transform 1 0 20064 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1036
timestamp 1626908933
transform 1 0 20064 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_232
timestamp 1626908933
transform 1 0 19488 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_830
timestamp 1626908933
transform 1 0 19488 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_635
timestamp 1626908933
transform 1 0 20832 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1626
timestamp 1626908933
transform 1 0 20832 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_16
timestamp 1626908933
transform 1 0 20832 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_78
timestamp 1626908933
transform 1 0 20832 0 -1 1332
box -38 -49 326 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_18
timestamp 1626908933
transform 1 0 20900 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_45
timestamp 1626908933
transform 1 0 20900 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_18
timestamp 1626908933
transform 1 0 20900 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_45
timestamp 1626908933
transform 1 0 20900 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_206
timestamp 1626908933
transform 1 0 20928 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_804
timestamp 1626908933
transform 1 0 20928 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_938
timestamp 1626908933
transform 1 0 21120 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_337
timestamp 1626908933
transform 1 0 21120 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1013
timestamp 1626908933
transform 1 0 21312 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1012
timestamp 1626908933
transform 1 0 21312 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_291
timestamp 1626908933
transform 1 0 21312 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_290
timestamp 1626908933
transform 1 0 21312 0 -1 1332
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_767
timestamp 1626908933
transform 1 0 22100 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_119
timestamp 1626908933
transform 1 0 22100 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_767
timestamp 1626908933
transform 1 0 22100 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_119
timestamp 1626908933
transform 1 0 22100 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_789
timestamp 1626908933
transform 1 0 22080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_788
timestamp 1626908933
transform 1 0 22080 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_191
timestamp 1626908933
transform 1 0 22080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_190
timestamp 1626908933
transform 1 0 22080 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_984
timestamp 1626908933
transform 1 0 22560 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_983
timestamp 1626908933
transform 1 0 22560 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_262
timestamp 1626908933
transform 1 0 22560 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_261
timestamp 1626908933
transform 1 0 22560 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_704
timestamp 1626908933
transform 1 0 22464 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_695
timestamp 1626908933
transform 1 0 22464 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_347
timestamp 1626908933
transform 1 0 22464 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_338
timestamp 1626908933
transform 1 0 22464 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_350
timestamp 1626908933
transform 1 0 23328 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_951
timestamp 1626908933
transform 1 0 23328 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_658
timestamp 1626908933
transform 1 0 23328 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1649
timestamp 1626908933
transform 1 0 23328 0 -1 1332
box -38 -49 134 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_17
timestamp 1626908933
transform 1 0 23300 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_44
timestamp 1626908933
transform 1 0 23300 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_17
timestamp 1626908933
transform 1 0 23300 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_44
timestamp 1626908933
transform 1 0 23300 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_12
timestamp 1626908933
transform 1 0 23424 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_73
timestamp 1626908933
transform 1 0 23424 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_336
timestamp 1626908933
transform 1 0 23712 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_937
timestamp 1626908933
transform 1 0 23712 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_165
timestamp 1626908933
transform 1 0 23520 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_763
timestamp 1626908933
transform 1 0 23520 0 1 0
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_743
timestamp 1626908933
transform 1 0 24500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_95
timestamp 1626908933
transform 1 0 24500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_743
timestamp 1626908933
transform 1 0 24500 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_95
timestamp 1626908933
transform 1 0 24500 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_951
timestamp 1626908933
transform 1 0 23904 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_950
timestamp 1626908933
transform 1 0 23904 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_229
timestamp 1626908933
transform 1 0 23904 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_228
timestamp 1626908933
transform 1 0 23904 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1643
timestamp 1626908933
transform 1 0 24864 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1609
timestamp 1626908933
transform 1 0 24672 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_652
timestamp 1626908933
transform 1 0 24864 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_618
timestamp 1626908933
transform 1 0 24672 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_950
timestamp 1626908933
transform 1 0 24672 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_349
timestamp 1626908933
transform 1 0 24672 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_738
timestamp 1626908933
transform 1 0 24768 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_140
timestamp 1626908933
transform 1 0 24768 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_346
timestamp 1626908933
transform 1 0 24960 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_703
timestamp 1626908933
transform 1 0 24960 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_634
timestamp 1626908933
transform 1 0 25056 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1625
timestamp 1626908933
transform 1 0 25056 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA2  fine_freq_track_VIA2_16
timestamp 1626908933
transform 1 0 25700 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_43
timestamp 1626908933
transform 1 0 25700 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_16
timestamp 1626908933
transform 1 0 25700 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_43
timestamp 1626908933
transform 1 0 25700 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_197
timestamp 1626908933
transform 1 0 25152 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_198
timestamp 1626908933
transform 1 0 25152 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_919
timestamp 1626908933
transform 1 0 25152 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_920
timestamp 1626908933
transform 1 0 25152 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_335
timestamp 1626908933
transform 1 0 25920 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_348
timestamp 1626908933
transform 1 0 25920 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_936
timestamp 1626908933
transform 1 0 25920 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_949
timestamp 1626908933
transform 1 0 25920 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_169
timestamp 1626908933
transform 1 0 26496 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_170
timestamp 1626908933
transform 1 0 26496 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_891
timestamp 1626908933
transform 1 0 26496 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_892
timestamp 1626908933
transform 1 0 26496 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_114
timestamp 1626908933
transform 1 0 26112 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_115
timestamp 1626908933
transform 1 0 26112 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_712
timestamp 1626908933
transform 1 0 26112 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_713
timestamp 1626908933
transform 1 0 26112 0 1 0
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_71
timestamp 1626908933
transform 1 0 26900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_719
timestamp 1626908933
transform 1 0 26900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_71
timestamp 1626908933
transform 1 0 26900 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_719
timestamp 1626908933
transform 1 0 26900 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_617
timestamp 1626908933
transform 1 0 27264 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_633
timestamp 1626908933
transform 1 0 27264 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_653
timestamp 1626908933
transform 1 0 27360 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_659
timestamp 1626908933
transform 1 0 27360 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1608
timestamp 1626908933
transform 1 0 27264 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1624
timestamp 1626908933
transform 1 0 27264 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1644
timestamp 1626908933
transform 1 0 27360 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1650
timestamp 1626908933
transform 1 0 27360 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_948
timestamp 1626908933
transform 1 0 27552 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_935
timestamp 1626908933
transform 1 0 27552 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_347
timestamp 1626908933
transform 1 0 27552 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_334
timestamp 1626908933
transform 1 0 27552 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_702
timestamp 1626908933
transform 1 0 27456 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_694
timestamp 1626908933
transform 1 0 27456 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_345
timestamp 1626908933
transform 1 0 27456 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_337
timestamp 1626908933
transform 1 0 27456 0 -1 1332
box -38 -49 134 715
use fine_freq_track_VIA3  fine_freq_track_VIA3_42
timestamp 1626908933
transform 1 0 28100 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_15
timestamp 1626908933
transform 1 0 28100 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_42
timestamp 1626908933
transform 1 0 28100 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_15
timestamp 1626908933
transform 1 0 28100 0 1 16
box -100 -33 100 33
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_861
timestamp 1626908933
transform 1 0 27744 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_860
timestamp 1626908933
transform 1 0 27744 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_139
timestamp 1626908933
transform 1 0 27744 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_138
timestamp 1626908933
transform 1 0 27744 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_616
timestamp 1626908933
transform 1 0 28896 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_632
timestamp 1626908933
transform 1 0 28896 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1607
timestamp 1626908933
transform 1 0 28896 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1623
timestamp 1626908933
transform 1 0 28896 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_47
timestamp 1626908933
transform 1 0 29300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_695
timestamp 1626908933
transform 1 0 29300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_47
timestamp 1626908933
transform 1 0 29300 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_695
timestamp 1626908933
transform 1 0 29300 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_103
timestamp 1626908933
transform 1 0 28992 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_104
timestamp 1626908933
transform 1 0 28992 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_825
timestamp 1626908933
transform 1 0 28992 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_826
timestamp 1626908933
transform 1 0 28992 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_70
timestamp 1626908933
transform 1 0 28512 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_71
timestamp 1626908933
transform 1 0 28512 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_668
timestamp 1626908933
transform 1 0 28512 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_669
timestamp 1626908933
transform 1 0 28512 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_333
timestamp 1626908933
transform 1 0 29760 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_934
timestamp 1626908933
transform 1 0 29760 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_631
timestamp 1626908933
transform 1 0 29760 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1622
timestamp 1626908933
transform 1 0 29760 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_344
timestamp 1626908933
transform 1 0 29952 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_701
timestamp 1626908933
transform 1 0 29952 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_346
timestamp 1626908933
transform 1 0 30048 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_947
timestamp 1626908933
transform 1 0 30048 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_654
timestamp 1626908933
transform 1 0 29856 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1645
timestamp 1626908933
transform 1 0 29856 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_38
timestamp 1626908933
transform 1 0 29952 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_636
timestamp 1626908933
transform 1 0 29952 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1621
timestamp 1626908933
transform 1 0 30240 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_630
timestamp 1626908933
transform 1 0 30240 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_790
timestamp 1626908933
transform 1 0 30336 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_789
timestamp 1626908933
transform 1 0 30336 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_68
timestamp 1626908933
transform 1 0 30336 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_67
timestamp 1626908933
transform 1 0 30336 0 -1 1332
box -38 -49 806 715
use fine_freq_track_VIA3  fine_freq_track_VIA3_41
timestamp 1626908933
transform 1 0 30500 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_14
timestamp 1626908933
transform 1 0 30500 0 1 23
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_41
timestamp 1626908933
transform 1 0 30500 0 1 16
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_14
timestamp 1626908933
transform 1 0 30500 0 1 16
box -100 -33 100 33
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_615
timestamp 1626908933
transform 1 0 31104 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_614
timestamp 1626908933
transform 1 0 31104 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_17
timestamp 1626908933
transform 1 0 31104 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_16
timestamp 1626908933
transform 1 0 31104 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_615
timestamp 1626908933
transform 1 0 31488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_629
timestamp 1626908933
transform 1 0 31488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1606
timestamp 1626908933
transform 1 0 31488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1620
timestamp 1626908933
transform 1 0 31488 0 1 0
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_671
timestamp 1626908933
transform 1 0 31700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_23
timestamp 1626908933
transform 1 0 31700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_671
timestamp 1626908933
transform 1 0 31700 0 1 666
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_23
timestamp 1626908933
transform 1 0 31700 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1651
timestamp 1626908933
transform 1 0 31584 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1646
timestamp 1626908933
transform 1 0 31584 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_660
timestamp 1626908933
transform 1 0 31584 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_655
timestamp 1626908933
transform 1 0 31584 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_700
timestamp 1626908933
transform 1 0 31680 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_693
timestamp 1626908933
transform 1 0 31680 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_343
timestamp 1626908933
transform 1 0 31680 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_336
timestamp 1626908933
transform 1 0 31680 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_357
timestamp 1626908933
transform 1 0 31776 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_359
timestamp 1626908933
transform 1 0 31776 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_958
timestamp 1626908933
transform 1 0 31776 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_960
timestamp 1626908933
transform 1 0 31776 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1652
timestamp 1626908933
transform 1 0 31968 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1647
timestamp 1626908933
transform 1 0 31968 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_661
timestamp 1626908933
transform 1 0 31968 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_656
timestamp 1626908933
transform 1 0 31968 0 1 0
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3929
timestamp 1626908933
transform 1 0 144 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1962
timestamp 1626908933
transform 1 0 144 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1653
timestamp 1626908933
transform 1 0 192 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_662
timestamp 1626908933
transform 1 0 192 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_692
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_335
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_961
timestamp 1626908933
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_360
timestamp 1626908933
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1192
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_594
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_698
timestamp 1626908933
transform 1 0 768 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1420
timestamp 1626908933
transform 1 0 768 0 1 1332
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1295
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_647
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1295
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_647
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1158
timestamp 1626908933
transform 1 0 1536 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_560
timestamp 1626908933
transform 1 0 1536 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_15
timestamp 1626908933
transform 1 0 2688 0 1 1332
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_7
timestamp 1626908933
transform 1 0 2688 0 1 1332
box -38 -49 902 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1386
timestamp 1626908933
transform 1 0 1920 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_664
timestamp 1626908933
transform 1 0 1920 0 1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3866
timestamp 1626908933
transform 1 0 3312 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2292
timestamp 1626908933
transform 1 0 3312 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1931
timestamp 1626908933
transform 1 0 3312 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_357
timestamp 1626908933
transform 1 0 3312 0 1 925
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2299
timestamp 1626908933
transform 1 0 3600 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_332
timestamp 1626908933
transform 1 0 3600 0 1 925
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1605
timestamp 1626908933
transform 1 0 3552 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_614
timestamp 1626908933
transform 1 0 3552 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1309
timestamp 1626908933
transform 1 0 3696 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3244
timestamp 1626908933
transform 1 0 3696 0 1 999
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_623
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1271
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_623
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1271
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_634
timestamp 1626908933
transform 1 0 4032 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1356
timestamp 1626908933
transform 1 0 4032 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_528
timestamp 1626908933
transform 1 0 3648 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1126
timestamp 1626908933
transform 1 0 3648 0 1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3716
timestamp 1626908933
transform 1 0 4560 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3243
timestamp 1626908933
transform 1 0 4464 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1781
timestamp 1626908933
transform 1 0 4560 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1308
timestamp 1626908933
transform 1 0 4464 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1604
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_613
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3237
timestamp 1626908933
transform 1 0 4848 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1302
timestamp 1626908933
transform 1 0 4848 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3192
timestamp 1626908933
transform 1 0 4848 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1225
timestamp 1626908933
transform 1 0 4848 0 1 1221
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_334
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_691
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_663
timestamp 1626908933
transform 1 0 4896 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1654
timestamp 1626908933
transform 1 0 4896 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1766
timestamp 1626908933
transform 1 0 4944 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3733
timestamp 1626908933
transform 1 0 4944 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_507
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1105
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_4
timestamp 1626908933
transform -1 0 5952 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_12
timestamp 1626908933
transform -1 0 5952 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_15
timestamp 1626908933
transform 1 0 5952 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_7
timestamp 1626908933
transform 1 0 5952 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_485
timestamp 1626908933
transform 1 0 6432 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1083
timestamp 1626908933
transform 1 0 6432 0 1 1332
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_599
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1247
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_599
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1247
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_664
timestamp 1626908933
transform 1 0 6816 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1655
timestamp 1626908933
transform 1 0 6816 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_27
timestamp 1626908933
transform 1 0 6912 0 1 1332
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_3
timestamp 1626908933
transform 1 0 6912 0 1 1332
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1223
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_575
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1223
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_575
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1251
timestamp 1626908933
transform 1 0 9216 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_529
timestamp 1626908933
transform 1 0 9216 0 1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2793
timestamp 1626908933
transform 1 0 10704 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_826
timestamp 1626908933
transform 1 0 10704 0 1 1073
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1656
timestamp 1626908933
transform 1 0 10080 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_665
timestamp 1626908933
transform 1 0 10080 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_690
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_333
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_29
timestamp 1626908933
transform 1 0 10176 0 1 1332
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_5
timestamp 1626908933
transform 1 0 10176 0 1 1332
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1199
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_551
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1199
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_551
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1979
timestamp 1626908933
transform 1 0 12432 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_44
timestamp 1626908933
transform 1 0 12432 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_972
timestamp 1626908933
transform 1 0 12480 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_374
timestamp 1626908933
transform 1 0 12480 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_612
timestamp 1626908933
transform 1 0 12864 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1603
timestamp 1626908933
transform 1 0 12864 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2802
timestamp 1626908933
transform 1 0 13296 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_867
timestamp 1626908933
transform 1 0 13296 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2790
timestamp 1626908933
transform 1 0 13200 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_823
timestamp 1626908933
transform 1 0 13200 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2796
timestamp 1626908933
transform 1 0 13200 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_861
timestamp 1626908933
transform 1 0 13200 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1977
timestamp 1626908933
transform 1 0 13488 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_42
timestamp 1626908933
transform 1 0 13488 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2007
timestamp 1626908933
transform 1 0 13488 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_40
timestamp 1626908933
transform 1 0 13488 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2006
timestamp 1626908933
transform 1 0 13488 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_39
timestamp 1626908933
transform 1 0 13488 0 1 1443
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_466
timestamp 1626908933
transform 1 0 12960 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1188
timestamp 1626908933
transform 1 0 12960 0 1 1332
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1175
timestamp 1626908933
transform 1 0 13700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_527
timestamp 1626908933
transform 1 0 13700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1175
timestamp 1626908933
transform 1 0 13700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_527
timestamp 1626908933
transform 1 0 13700 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_933
timestamp 1626908933
transform 1 0 13728 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_332
timestamp 1626908933
transform 1 0 13728 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_361
timestamp 1626908933
transform 1 0 14016 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_962
timestamp 1626908933
transform 1 0 14016 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_611
timestamp 1626908933
transform 1 0 13920 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_666
timestamp 1626908933
transform 1 0 14208 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1602
timestamp 1626908933
transform 1 0 13920 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1657
timestamp 1626908933
transform 1 0 14208 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_828
timestamp 1626908933
transform 1 0 14640 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2795
timestamp 1626908933
transform 1 0 14640 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_40
timestamp 1626908933
transform 1 0 14256 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1975
timestamp 1626908933
transform 1 0 14256 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_2
timestamp 1626908933
transform -1 0 14880 0 1 1332
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_41
timestamp 1626908933
transform -1 0 14880 0 1 1332
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1658
timestamp 1626908933
transform 1 0 14880 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1601
timestamp 1626908933
transform 1 0 15456 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_667
timestamp 1626908933
transform 1 0 14880 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_610
timestamp 1626908933
transform 1 0 15456 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_923
timestamp 1626908933
transform 1 0 15072 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_325
timestamp 1626908933
transform 1 0 15072 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_689
timestamp 1626908933
transform 1 0 14976 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_332
timestamp 1626908933
transform 1 0 14976 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_831
timestamp 1626908933
transform 1 0 15600 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2798
timestamp 1626908933
transform 1 0 15600 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_865
timestamp 1626908933
transform 1 0 15792 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_871
timestamp 1626908933
transform 1 0 15888 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2800
timestamp 1626908933
transform 1 0 15792 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2806
timestamp 1626908933
transform 1 0 15888 0 1 1221
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_609
timestamp 1626908933
transform 1 0 16320 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1600
timestamp 1626908933
transform 1 0 16320 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_742
timestamp 1626908933
transform 1 0 15984 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2677
timestamp 1626908933
transform 1 0 15984 0 1 999
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_503
timestamp 1626908933
transform 1 0 16100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1151
timestamp 1626908933
transform 1 0 16100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_503
timestamp 1626908933
transform 1 0 16100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1151
timestamp 1626908933
transform 1 0 16100 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_417
timestamp 1626908933
transform 1 0 15552 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1139
timestamp 1626908933
transform 1 0 15552 0 1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2685
timestamp 1626908933
transform 1 0 16464 0 1 1147
box -32 -32 32 32
use M1M2_PR  M1M2_PR_718
timestamp 1626908933
transform 1 0 16464 0 1 1147
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_896
timestamp 1626908933
transform 1 0 16416 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_298
timestamp 1626908933
transform 1 0 16416 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1109
timestamp 1626908933
transform 1 0 16800 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_387
timestamp 1626908933
transform 1 0 16800 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_608
timestamp 1626908933
transform 1 0 17568 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1599
timestamp 1626908933
transform 1 0 17568 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2799
timestamp 1626908933
transform 1 0 17904 0 1 851
box -29 -23 29 23
use L1M1_PR  L1M1_PR_864
timestamp 1626908933
transform 1 0 17904 0 1 851
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3490
timestamp 1626908933
transform 1 0 18192 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2674
timestamp 1626908933
transform 1 0 18096 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1555
timestamp 1626908933
transform 1 0 18192 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_739
timestamp 1626908933
transform 1 0 18096 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3438
timestamp 1626908933
transform 1 0 18192 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1471
timestamp 1626908933
transform 1 0 18192 0 1 1221
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1598
timestamp 1626908933
transform 1 0 18048 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_607
timestamp 1626908933
transform 1 0 18048 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_364
timestamp 1626908933
transform 1 0 18144 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1086
timestamp 1626908933
transform 1 0 18144 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_276
timestamp 1626908933
transform 1 0 17664 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_874
timestamp 1626908933
transform 1 0 17664 0 1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_868
timestamp 1626908933
transform 1 0 18288 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2803
timestamp 1626908933
transform 1 0 18288 0 1 1073
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_479
timestamp 1626908933
transform 1 0 18500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1127
timestamp 1626908933
transform 1 0 18500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_479
timestamp 1626908933
transform 1 0 18500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1127
timestamp 1626908933
transform 1 0 18500 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_331
timestamp 1626908933
transform 1 0 18912 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_932
timestamp 1626908933
transform 1 0 18912 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_606
timestamp 1626908933
transform 1 0 19104 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1597
timestamp 1626908933
transform 1 0 19104 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1055
timestamp 1626908933
transform 1 0 19200 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_333
timestamp 1626908933
transform 1 0 19200 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1034
timestamp 1626908933
transform 1 0 20064 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_312
timestamp 1626908933
transform 1 0 20064 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_688
timestamp 1626908933
transform 1 0 19968 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_331
timestamp 1626908933
transform 1 0 19968 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_739
timestamp 1626908933
transform 1 0 20976 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2706
timestamp 1626908933
transform 1 0 20976 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_762
timestamp 1626908933
transform 1 0 20880 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2697
timestamp 1626908933
transform 1 0 20880 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_894
timestamp 1626908933
transform 1 0 20688 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2861
timestamp 1626908933
transform 1 0 20688 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_940
timestamp 1626908933
transform 1 0 20976 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2875
timestamp 1626908933
transform 1 0 20976 0 1 1221
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_455
timestamp 1626908933
transform 1 0 20900 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1103
timestamp 1626908933
transform 1 0 20900 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_455
timestamp 1626908933
transform 1 0 20900 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1103
timestamp 1626908933
transform 1 0 20900 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_24
timestamp 1626908933
transform -1 0 21216 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_86
timestamp 1626908933
transform -1 0 21216 0 1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2874
timestamp 1626908933
transform 1 0 21072 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_939
timestamp 1626908933
transform 1 0 21072 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2857
timestamp 1626908933
transform 1 0 21264 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_890
timestamp 1626908933
transform 1 0 21264 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1596
timestamp 1626908933
transform 1 0 21216 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_605
timestamp 1626908933
transform 1 0 21216 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1011
timestamp 1626908933
transform 1 0 21312 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_289
timestamp 1626908933
transform 1 0 21312 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_787
timestamp 1626908933
transform 1 0 22080 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_189
timestamp 1626908933
transform 1 0 22080 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1595
timestamp 1626908933
transform 1 0 22464 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_604
timestamp 1626908933
transform 1 0 22464 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_982
timestamp 1626908933
transform 1 0 22560 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_260
timestamp 1626908933
transform 1 0 22560 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_603
timestamp 1626908933
transform 1 0 23328 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1594
timestamp 1626908933
transform 1 0 23328 0 1 1332
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_431
timestamp 1626908933
transform 1 0 23300 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1079
timestamp 1626908933
transform 1 0 23300 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_431
timestamp 1626908933
transform 1 0 23300 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1079
timestamp 1626908933
transform 1 0 23300 0 1 1332
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2869
timestamp 1626908933
transform 1 0 23472 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_934
timestamp 1626908933
transform 1 0 23472 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2853
timestamp 1626908933
transform 1 0 23472 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_886
timestamp 1626908933
transform 1 0 23472 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2872
timestamp 1626908933
transform 1 0 23568 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2051
timestamp 1626908933
transform 1 0 23664 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_937
timestamp 1626908933
transform 1 0 23568 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_116
timestamp 1626908933
transform 1 0 23664 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2070
timestamp 1626908933
transform 1 0 23664 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_103
timestamp 1626908933
transform 1 0 23664 0 1 1073
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_164
timestamp 1626908933
transform 1 0 23424 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_762
timestamp 1626908933
transform 1 0 23424 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_10
timestamp 1626908933
transform -1 0 24384 0 1 1332
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_49
timestamp 1626908933
transform -1 0 24384 0 1 1332
box -38 -49 614 715
use M1M2_PR  M1M2_PR_2855
timestamp 1626908933
transform 1 0 24144 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_888
timestamp 1626908933
transform 1 0 24144 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_742
timestamp 1626908933
transform 1 0 24384 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_144
timestamp 1626908933
transform 1 0 24384 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_963
timestamp 1626908933
transform 1 0 24768 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_362
timestamp 1626908933
transform 1 0 24768 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_330
timestamp 1626908933
transform 1 0 24960 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_687
timestamp 1626908933
transform 1 0 24960 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_602
timestamp 1626908933
transform 1 0 25056 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1593
timestamp 1626908933
transform 1 0 25056 0 1 1332
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_407
timestamp 1626908933
transform 1 0 25700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1055
timestamp 1626908933
transform 1 0 25700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_407
timestamp 1626908933
transform 1 0 25700 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1055
timestamp 1626908933
transform 1 0 25700 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_196
timestamp 1626908933
transform 1 0 25152 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_918
timestamp 1626908933
transform 1 0 25152 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_931
timestamp 1626908933
transform 1 0 25920 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_330
timestamp 1626908933
transform 1 0 25920 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_711
timestamp 1626908933
transform 1 0 26112 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_113
timestamp 1626908933
transform 1 0 26112 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_890
timestamp 1626908933
transform 1 0 26496 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_168
timestamp 1626908933
transform 1 0 26496 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1592
timestamp 1626908933
transform 1 0 27264 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_601
timestamp 1626908933
transform 1 0 27264 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_687
timestamp 1626908933
transform 1 0 27360 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_89
timestamp 1626908933
transform 1 0 27360 0 1 1332
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1031
timestamp 1626908933
transform 1 0 28100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_383
timestamp 1626908933
transform 1 0 28100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1031
timestamp 1626908933
transform 1 0 28100 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_383
timestamp 1626908933
transform 1 0 28100 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_859
timestamp 1626908933
transform 1 0 27744 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_137
timestamp 1626908933
transform 1 0 27744 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1591
timestamp 1626908933
transform 1 0 28896 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_600
timestamp 1626908933
transform 1 0 28896 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_667
timestamp 1626908933
transform 1 0 28512 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_69
timestamp 1626908933
transform 1 0 28512 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_824
timestamp 1626908933
transform 1 0 28992 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_102
timestamp 1626908933
transform 1 0 28992 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1659
timestamp 1626908933
transform 1 0 29856 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1590
timestamp 1626908933
transform 1 0 29760 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_668
timestamp 1626908933
transform 1 0 29856 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_599
timestamp 1626908933
transform 1 0 29760 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_930
timestamp 1626908933
transform 1 0 30048 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_329
timestamp 1626908933
transform 1 0 30048 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_686
timestamp 1626908933
transform 1 0 29952 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_329
timestamp 1626908933
transform 1 0 29952 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1589
timestamp 1626908933
transform 1 0 30240 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_598
timestamp 1626908933
transform 1 0 30240 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_788
timestamp 1626908933
transform 1 0 30336 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_66
timestamp 1626908933
transform 1 0 30336 0 1 1332
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1007
timestamp 1626908933
transform 1 0 30500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_359
timestamp 1626908933
transform 1 0 30500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1007
timestamp 1626908933
transform 1 0 30500 0 1 1332
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_359
timestamp 1626908933
transform 1 0 30500 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1588
timestamp 1626908933
transform 1 0 31104 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_597
timestamp 1626908933
transform 1 0 31104 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_744
timestamp 1626908933
transform 1 0 31200 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_22
timestamp 1626908933
transform 1 0 31200 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1660
timestamp 1626908933
transform 1 0 31968 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_669
timestamp 1626908933
transform 1 0 31968 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_328
timestamp 1626908933
transform 1 0 0 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_929
timestamp 1626908933
transform 1 0 0 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1961
timestamp 1626908933
transform 1 0 48 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3928
timestamp 1626908933
transform 1 0 48 0 1 1665
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_334
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_982
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_334
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_982
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_720
timestamp 1626908933
transform 1 0 192 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1442
timestamp 1626908933
transform 1 0 192 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1587
timestamp 1626908933
transform 1 0 960 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_596
timestamp 1626908933
transform 1 0 960 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1181
timestamp 1626908933
transform 1 0 1056 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_583
timestamp 1626908933
transform 1 0 1056 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1409
timestamp 1626908933
transform 1 0 1440 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_687
timestamp 1626908933
transform 1 0 1440 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1586
timestamp 1626908933
transform 1 0 2208 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_595
timestamp 1626908933
transform 1 0 2208 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_964
timestamp 1626908933
transform 1 0 2304 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_363
timestamp 1626908933
transform 1 0 2304 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_685
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_328
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3927
timestamp 1626908933
transform 1 0 2736 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3926
timestamp 1626908933
transform 1 0 2736 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1960
timestamp 1626908933
transform 1 0 2736 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1959
timestamp 1626908933
transform 1 0 2736 0 1 2257
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_965
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_364
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_958
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_310
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_958
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_310
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3865
timestamp 1626908933
transform 1 0 2832 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1930
timestamp 1626908933
transform 1 0 2832 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1661
timestamp 1626908933
transform 1 0 2784 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_670
timestamp 1626908933
transform 1 0 2784 0 -1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3864
timestamp 1626908933
transform 1 0 3120 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1929
timestamp 1626908933
transform 1 0 3120 0 1 2257
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3717
timestamp 1626908933
transform 1 0 3120 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1750
timestamp 1626908933
transform 1 0 3120 0 1 1887
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3695
timestamp 1626908933
transform 1 0 3216 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3290
timestamp 1626908933
transform 1 0 3312 0 1 2183
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1760
timestamp 1626908933
transform 1 0 3216 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1355
timestamp 1626908933
transform 1 0 3312 0 1 2183
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_594
timestamp 1626908933
transform 1 0 3552 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1585
timestamp 1626908933
transform 1 0 3552 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_329
timestamp 1626908933
transform 1 0 3408 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1268
timestamp 1626908933
transform 1 0 3504 0 1 2183
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2296
timestamp 1626908933
transform 1 0 3408 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3235
timestamp 1626908933
transform 1 0 3504 0 1 2183
box -32 -32 32 32
use L1M1_PR  L1M1_PR_354
timestamp 1626908933
transform 1 0 3408 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2289
timestamp 1626908933
transform 1 0 3408 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__o21ai_2  sky130_fd_sc_hs__o21ai_2_0
timestamp 1626908933
transform -1 0 3552 0 -1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__o21ai_2  sky130_fd_sc_hs__o21ai_2_1
timestamp 1626908933
transform -1 0 3552 0 -1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_633
timestamp 1626908933
transform 1 0 3648 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1355
timestamp 1626908933
transform 1 0 3648 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__nand2b_4  sky130_fd_sc_hs__nand2b_4_1
timestamp 1626908933
transform 1 0 4416 0 -1 2664
box -38 -49 1190 715
use sky130_fd_sc_hs__nand2b_4  sky130_fd_sc_hs__nand2b_4_0
timestamp 1626908933
transform 1 0 4416 0 -1 2664
box -38 -49 1190 715
use L1M1_PR  L1M1_PR_3715
timestamp 1626908933
transform 1 0 4944 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1780
timestamp 1626908933
transform 1 0 4944 0 1 2109
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3924
timestamp 1626908933
transform 1 0 4560 0 1 1739
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3732
timestamp 1626908933
transform 1 0 4944 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1957
timestamp 1626908933
transform 1 0 4560 0 1 1739
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1765
timestamp 1626908933
transform 1 0 4944 0 1 2109
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_934
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_286
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_934
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_286
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2360
timestamp 1626908933
transform 1 0 5616 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_425
timestamp 1626908933
transform 1 0 5616 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3861
timestamp 1626908933
transform 1 0 5808 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3260
timestamp 1626908933
transform 1 0 5808 0 1 1813
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1926
timestamp 1626908933
transform 1 0 5808 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1325
timestamp 1626908933
transform 1 0 5808 0 1 1813
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1662
timestamp 1626908933
transform 1 0 5760 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_671
timestamp 1626908933
transform 1 0 5760 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_966
timestamp 1626908933
transform 1 0 5568 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_365
timestamp 1626908933
transform 1 0 5568 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_427
timestamp 1626908933
transform 1 0 6000 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2394
timestamp 1626908933
transform 1 0 6000 0 1 1591
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1924
timestamp 1626908933
transform 1 0 6096 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3859
timestamp 1626908933
transform 1 0 6096 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_423
timestamp 1626908933
transform 1 0 6288 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2358
timestamp 1626908933
transform 1 0 6288 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1758
timestamp 1626908933
transform 1 0 6192 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3725
timestamp 1626908933
transform 1 0 6192 0 1 1887
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1769
timestamp 1626908933
transform 1 0 6096 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3704
timestamp 1626908933
transform 1 0 6096 0 1 1887
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_928
timestamp 1626908933
transform 1 0 6336 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_327
timestamp 1626908933
transform 1 0 6336 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_5
timestamp 1626908933
transform 1 0 5856 0 -1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_11
timestamp 1626908933
transform 1 0 5856 0 -1 2664
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1242
timestamp 1626908933
transform 1 0 6672 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1475
timestamp 1626908933
transform 1 0 7056 0 1 1739
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3209
timestamp 1626908933
transform 1 0 6672 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3442
timestamp 1626908933
transform 1 0 7056 0 1 1739
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1562
timestamp 1626908933
transform 1 0 6960 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3497
timestamp 1626908933
transform 1 0 6960 0 1 1739
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1474
timestamp 1626908933
transform 1 0 7056 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3441
timestamp 1626908933
transform 1 0 7056 0 1 2109
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_583
timestamp 1626908933
transform 1 0 6528 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1305
timestamp 1626908933
transform 1 0 6528 0 -1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3849
timestamp 1626908933
transform 1 0 7344 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1914
timestamp 1626908933
transform 1 0 7344 0 1 1665
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_910
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_262
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_910
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_262
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_684
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_327
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_927
timestamp 1626908933
transform 1 0 7296 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_326
timestamp 1626908933
transform 1 0 7296 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1943
timestamp 1626908933
transform 1 0 7920 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3910
timestamp 1626908933
transform 1 0 7920 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_561
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1283
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_819
timestamp 1626908933
transform 1 0 8688 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2786
timestamp 1626908933
transform 1 0 8688 0 1 2257
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1561
timestamp 1626908933
transform 1 0 8400 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3496
timestamp 1626908933
transform 1 0 8400 0 1 2109
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_325
timestamp 1626908933
transform 1 0 8928 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_926
timestamp 1626908933
transform 1 0 8928 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_33
timestamp 1626908933
transform 1 0 8880 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2000
timestamp 1626908933
transform 1 0 8880 0 1 1887
box -32 -32 32 32
use L1M1_PR  L1M1_PR_854
timestamp 1626908933
transform 1 0 8784 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2789
timestamp 1626908933
transform 1 0 8784 0 1 2257
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_541
timestamp 1626908933
transform 1 0 9120 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1263
timestamp 1626908933
transform 1 0 9120 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_1
timestamp 1626908933
transform 1 0 8352 0 -1 2664
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_40
timestamp 1626908933
transform 1 0 8352 0 -1 2664
box -38 -49 614 715
use L1M1_PR  L1M1_PR_1969
timestamp 1626908933
transform 1 0 9168 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_34
timestamp 1626908933
transform 1 0 9168 0 1 1887
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_60
timestamp 1626908933
transform 1 0 9888 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_8
timestamp 1626908933
transform 1 0 9888 0 -1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3493
timestamp 1626908933
transform 1 0 10224 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1558
timestamp 1626908933
transform 1 0 10224 0 1 1591
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3695
timestamp 1626908933
transform 1 0 10320 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1728
timestamp 1626908933
transform 1 0 10320 0 1 1813
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_886
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_238
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_886
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_238
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_925
timestamp 1626908933
transform 1 0 10272 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_324
timestamp 1626908933
transform 1 0 10272 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_672
timestamp 1626908933
transform 1 0 10464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1663
timestamp 1626908933
transform 1 0 10464 0 -1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1907
timestamp 1626908933
transform 1 0 10608 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3842
timestamp 1626908933
transform 1 0 10608 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_25
timestamp 1626908933
transform -1 0 10848 0 -1 2664
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_87
timestamp 1626908933
transform -1 0 10848 0 -1 2664
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_924
timestamp 1626908933
transform 1 0 10848 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_323
timestamp 1626908933
transform 1 0 10848 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1221
timestamp 1626908933
transform 1 0 11040 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_499
timestamp 1626908933
transform 1 0 11040 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_322
timestamp 1626908933
transform 1 0 11808 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_923
timestamp 1626908933
transform 1 0 11808 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_383
timestamp 1626908933
transform 1 0 12096 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_981
timestamp 1626908933
transform 1 0 12096 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_593
timestamp 1626908933
transform 1 0 12000 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1584
timestamp 1626908933
transform 1 0 12000 0 -1 2664
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_214
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_862
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_214
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_862
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2789
timestamp 1626908933
transform 1 0 13200 0 1 1739
box -32 -32 32 32
use M1M2_PR  M1M2_PR_822
timestamp 1626908933
transform 1 0 13200 0 1 1739
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1664
timestamp 1626908933
transform 1 0 12576 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_673
timestamp 1626908933
transform 1 0 12576 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_683
timestamp 1626908933
transform 1 0 12480 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_326
timestamp 1626908933
transform 1 0 12480 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_30
timestamp 1626908933
transform -1 0 14880 0 -1 2664
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_5
timestamp 1626908933
transform -1 0 14880 0 -1 2664
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_860
timestamp 1626908933
transform 1 0 14448 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2795
timestamp 1626908933
transform 1 0 14448 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3492
timestamp 1626908933
transform 1 0 14832 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2801
timestamp 1626908933
transform 1 0 14640 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1557
timestamp 1626908933
transform 1 0 14832 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_866
timestamp 1626908933
transform 1 0 14640 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2794
timestamp 1626908933
transform 1 0 14640 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_827
timestamp 1626908933
transform 1 0 14640 0 1 1665
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_838
timestamp 1626908933
transform 1 0 14900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_190
timestamp 1626908933
transform 1 0 14900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_838
timestamp 1626908933
transform 1 0 14900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_190
timestamp 1626908933
transform 1 0 14900 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_967
timestamp 1626908933
transform 1 0 14880 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_366
timestamp 1626908933
transform 1 0 14880 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_674
timestamp 1626908933
transform 1 0 15072 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1665
timestamp 1626908933
transform 1 0 15072 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_30
timestamp 1626908933
transform -1 0 17472 0 -1 2664
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_6
timestamp 1626908933
transform -1 0 17472 0 -1 2664
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_814
timestamp 1626908933
transform 1 0 17300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_166
timestamp 1626908933
transform 1 0 17300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_814
timestamp 1626908933
transform 1 0 17300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_166
timestamp 1626908933
transform 1 0 17300 0 1 1998
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3491
timestamp 1626908933
transform 1 0 17424 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1556
timestamp 1626908933
transform 1 0 17424 0 1 2257
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_325
timestamp 1626908933
transform 1 0 17472 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_682
timestamp 1626908933
transform 1 0 17472 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_592
timestamp 1626908933
transform 1 0 17568 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1583
timestamp 1626908933
transform 1 0 17568 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_591
timestamp 1626908933
transform 1 0 18048 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1582
timestamp 1626908933
transform 1 0 18048 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1470
timestamp 1626908933
transform 1 0 18192 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3437
timestamp 1626908933
transform 1 0 18192 0 1 2257
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_363
timestamp 1626908933
transform 1 0 18144 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1085
timestamp 1626908933
transform 1 0 18144 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_275
timestamp 1626908933
transform 1 0 17664 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_873
timestamp 1626908933
transform 1 0 17664 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1581
timestamp 1626908933
transform 1 0 19104 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_590
timestamp 1626908933
transform 1 0 19104 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_922
timestamp 1626908933
transform 1 0 18912 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_321
timestamp 1626908933
transform 1 0 18912 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1054
timestamp 1626908933
transform 1 0 19200 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_332
timestamp 1626908933
transform 1 0 19200 0 -1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1439
timestamp 1626908933
transform 1 0 20112 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3406
timestamp 1626908933
transform 1 0 20112 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_893
timestamp 1626908933
transform 1 0 20688 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2860
timestamp 1626908933
transform 1 0 20688 0 1 1813
box -32 -32 32 32
use L1M1_PR  L1M1_PR_941
timestamp 1626908933
transform 1 0 20784 0 1 1813
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2876
timestamp 1626908933
transform 1 0 20784 0 1 1813
box -29 -23 29 23
use M1M2_PR  M1M2_PR_737
timestamp 1626908933
transform 1 0 21072 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2704
timestamp 1626908933
transform 1 0 21072 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_760
timestamp 1626908933
transform 1 0 21072 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2695
timestamp 1626908933
transform 1 0 21072 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_889
timestamp 1626908933
transform 1 0 21264 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2856
timestamp 1626908933
transform 1 0 21264 0 1 1591
box -32 -32 32 32
use L1M1_PR  L1M1_PR_938
timestamp 1626908933
transform 1 0 21168 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2873
timestamp 1626908933
transform 1 0 21168 0 1 1591
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_142
timestamp 1626908933
transform 1 0 19700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_790
timestamp 1626908933
transform 1 0 19700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_142
timestamp 1626908933
transform 1 0 19700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_790
timestamp 1626908933
transform 1 0 19700 0 1 1998
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1438
timestamp 1626908933
transform 1 0 20112 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3405
timestamp 1626908933
transform 1 0 20112 0 1 2257
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1524
timestamp 1626908933
transform 1 0 20016 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3459
timestamp 1626908933
transform 1 0 20016 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1523
timestamp 1626908933
transform 1 0 20880 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3458
timestamp 1626908933
transform 1 0 20880 0 1 1887
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_118
timestamp 1626908933
transform 1 0 22100 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_766
timestamp 1626908933
transform 1 0 22100 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_118
timestamp 1626908933
transform 1 0 22100 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_766
timestamp 1626908933
transform 1 0 22100 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_45
timestamp 1626908933
transform 1 0 19968 0 -1 2664
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_21
timestamp 1626908933
transform 1 0 19968 0 -1 2664
box -38 -49 2342 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_968
timestamp 1626908933
transform 1 0 22272 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_367
timestamp 1626908933
transform 1 0 22272 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_981
timestamp 1626908933
transform 1 0 22560 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_259
timestamp 1626908933
transform 1 0 22560 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_681
timestamp 1626908933
transform 1 0 22464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_324
timestamp 1626908933
transform 1 0 22464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_320
timestamp 1626908933
transform 1 0 23328 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_921
timestamp 1626908933
transform 1 0 23328 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_99
timestamp 1626908933
transform 1 0 23760 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_102
timestamp 1626908933
transform 1 0 23664 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_885
timestamp 1626908933
transform 1 0 23472 0 1 1739
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2066
timestamp 1626908933
transform 1 0 23760 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2069
timestamp 1626908933
transform 1 0 23664 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2852
timestamp 1626908933
transform 1 0 23472 0 1 1739
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_163
timestamp 1626908933
transform 1 0 23520 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_761
timestamp 1626908933
transform 1 0 23520 0 -1 2664
box -38 -49 422 715
use M1M2_PR  M1M2_PR_887
timestamp 1626908933
transform 1 0 24144 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2854
timestamp 1626908933
transform 1 0 24144 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_115
timestamp 1626908933
transform 1 0 23856 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_933
timestamp 1626908933
transform 1 0 23952 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_936
timestamp 1626908933
transform 1 0 24144 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2050
timestamp 1626908933
transform 1 0 23856 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2868
timestamp 1626908933
transform 1 0 23952 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2871
timestamp 1626908933
transform 1 0 24144 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1526
timestamp 1626908933
transform 1 0 24336 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3461
timestamp 1626908933
transform 1 0 24336 0 1 1887
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_94
timestamp 1626908933
transform 1 0 24500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_742
timestamp 1626908933
transform 1 0 24500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_94
timestamp 1626908933
transform 1 0 24500 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_742
timestamp 1626908933
transform 1 0 24500 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_227
timestamp 1626908933
transform 1 0 23904 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_949
timestamp 1626908933
transform 1 0 23904 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1666
timestamp 1626908933
transform 1 0 24864 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_675
timestamp 1626908933
transform 1 0 24864 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_920
timestamp 1626908933
transform 1 0 24672 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_319
timestamp 1626908933
transform 1 0 24672 0 -1 2664
box -38 -49 230 715
use L1M1_PR  L1M1_PR_2047
timestamp 1626908933
transform 1 0 25008 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_112
timestamp 1626908933
transform 1 0 25008 0 1 2109
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1685
timestamp 1626908933
transform 1 0 27024 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3652
timestamp 1626908933
transform 1 0 27024 0 1 2257
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_70
timestamp 1626908933
transform 1 0 26900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_718
timestamp 1626908933
transform 1 0 26900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_70
timestamp 1626908933
transform 1 0 26900 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_718
timestamp 1626908933
transform 1 0 26900 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_368
timestamp 1626908933
transform 1 0 27264 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_969
timestamp 1626908933
transform 1 0 27264 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1440
timestamp 1626908933
transform 1 0 27120 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1441
timestamp 1626908933
transform 1 0 27120 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3407
timestamp 1626908933
transform 1 0 27120 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3408
timestamp 1626908933
transform 1 0 27120 0 1 1887
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1525
timestamp 1626908933
transform 1 0 27216 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3460
timestamp 1626908933
transform 1 0 27216 0 1 2257
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_323
timestamp 1626908933
transform 1 0 27456 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_680
timestamp 1626908933
transform 1 0 27456 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_318
timestamp 1626908933
transform 1 0 27552 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_919
timestamp 1626908933
transform 1 0 27552 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_44
timestamp 1626908933
transform -1 0 27264 0 -1 2664
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_20
timestamp 1626908933
transform -1 0 27264 0 -1 2664
box -38 -49 2342 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_858
timestamp 1626908933
transform 1 0 27744 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_136
timestamp 1626908933
transform 1 0 27744 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_589
timestamp 1626908933
transform 1 0 28896 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1580
timestamp 1626908933
transform 1 0 28896 0 -1 2664
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_46
timestamp 1626908933
transform 1 0 29300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_694
timestamp 1626908933
transform 1 0 29300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_46
timestamp 1626908933
transform 1 0 29300 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_694
timestamp 1626908933
transform 1 0 29300 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_101
timestamp 1626908933
transform 1 0 28992 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_823
timestamp 1626908933
transform 1 0 28992 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_68
timestamp 1626908933
transform 1 0 28512 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_666
timestamp 1626908933
transform 1 0 28512 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_918
timestamp 1626908933
transform 1 0 29760 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_317
timestamp 1626908933
transform 1 0 29760 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_635
timestamp 1626908933
transform 1 0 29952 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_37
timestamp 1626908933
transform 1 0 29952 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_787
timestamp 1626908933
transform 1 0 30336 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_65
timestamp 1626908933
transform 1 0 30336 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_613
timestamp 1626908933
transform 1 0 31104 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_15
timestamp 1626908933
transform 1 0 31104 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_588
timestamp 1626908933
transform 1 0 31488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1579
timestamp 1626908933
transform 1 0 31488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_322
timestamp 1626908933
transform 1 0 31680 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_679
timestamp 1626908933
transform 1 0 31680 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_676
timestamp 1626908933
transform 1 0 31584 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1667
timestamp 1626908933
transform 1 0 31584 0 -1 2664
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_22
timestamp 1626908933
transform 1 0 31700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_670
timestamp 1626908933
transform 1 0 31700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_22
timestamp 1626908933
transform 1 0 31700 0 1 1998
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_670
timestamp 1626908933
transform 1 0 31700 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_369
timestamp 1626908933
transform 1 0 31776 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_970
timestamp 1626908933
transform 1 0 31776 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1668
timestamp 1626908933
transform 1 0 31968 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_677
timestamp 1626908933
transform 1 0 31968 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_321
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_678
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_370
timestamp 1626908933
transform 1 0 0 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_971
timestamp 1626908933
transform 1 0 0 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_678
timestamp 1626908933
transform 1 0 192 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1669
timestamp 1626908933
transform 1 0 192 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_697
timestamp 1626908933
transform 1 0 768 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1419
timestamp 1626908933
transform 1 0 768 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_593
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1191
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1294
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_646
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1294
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_646
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1578
timestamp 1626908933
transform 1 0 1536 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_587
timestamp 1626908933
transform 1 0 1536 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1157
timestamp 1626908933
transform 1 0 1632 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_559
timestamp 1626908933
transform 1 0 1632 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1577
timestamp 1626908933
transform 1 0 2016 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_586
timestamp 1626908933
transform 1 0 2016 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1385
timestamp 1626908933
transform 1 0 2112 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_663
timestamp 1626908933
transform 1 0 2112 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_585
timestamp 1626908933
transform 1 0 2880 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1576
timestamp 1626908933
transform 1 0 2880 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1238
timestamp 1626908933
transform 1 0 3120 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1749
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3205
timestamp 1626908933
transform 1 0 3120 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3716
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1761
timestamp 1626908933
transform 1 0 2928 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3696
timestamp 1626908933
transform 1 0 2928 0 1 2405
box -29 -23 29 23
use M1M2_PR  M1M2_PR_328
timestamp 1626908933
transform 1 0 3408 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1267
timestamp 1626908933
transform 1 0 3504 0 1 2849
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2295
timestamp 1626908933
transform 1 0 3408 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3234
timestamp 1626908933
transform 1 0 3504 0 1 2849
box -32 -32 32 32
use L1M1_PR  L1M1_PR_355
timestamp 1626908933
transform 1 0 3312 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2290
timestamp 1626908933
transform 1 0 3312 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_650
timestamp 1626908933
transform 1 0 3360 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1372
timestamp 1626908933
transform 1 0 3360 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_544
timestamp 1626908933
transform 1 0 2976 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1142
timestamp 1626908933
transform 1 0 2976 0 1 2664
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1270
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_622
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1270
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_622
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3256
timestamp 1626908933
transform 1 0 4272 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1321
timestamp 1626908933
transform 1 0 4272 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_3
timestamp 1626908933
transform 1 0 4128 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_11
timestamp 1626908933
transform 1 0 4128 0 1 2664
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1956
timestamp 1626908933
transform 1 0 4560 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3923
timestamp 1626908933
transform 1 0 4560 0 1 2405
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1319
timestamp 1626908933
transform 1 0 4464 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1928
timestamp 1626908933
transform 1 0 4464 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3254
timestamp 1626908933
transform 1 0 4464 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3863
timestamp 1626908933
transform 1 0 4464 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_320
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_677
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_371
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_972
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_679
timestamp 1626908933
transform 1 0 5280 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1670
timestamp 1626908933
transform 1 0 5280 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_522
timestamp 1626908933
transform 1 0 4608 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1120
timestamp 1626908933
transform 1 0 4608 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_120
timestamp 1626908933
transform 1 0 5376 0 1 2664
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_59
timestamp 1626908933
transform 1 0 5376 0 1 2664
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3288
timestamp 1626908933
transform 1 0 5616 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3287
timestamp 1626908933
transform 1 0 5616 0 1 2849
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2288
timestamp 1626908933
transform 1 0 5616 0 1 2479
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1353
timestamp 1626908933
transform 1 0 5616 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1352
timestamp 1626908933
transform 1 0 5616 0 1 2849
box -29 -23 29 23
use L1M1_PR  L1M1_PR_353
timestamp 1626908933
transform 1 0 5616 0 1 2479
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1575
timestamp 1626908933
transform 1 0 5664 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_584
timestamp 1626908933
transform 1 0 5664 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3860
timestamp 1626908933
transform 1 0 5904 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1925
timestamp 1626908933
transform 1 0 5904 0 1 2405
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2294
timestamp 1626908933
transform 1 0 5904 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_327
timestamp 1626908933
transform 1 0 5904 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2393
timestamp 1626908933
transform 1 0 6000 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_426
timestamp 1626908933
transform 1 0 6000 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3703
timestamp 1626908933
transform 1 0 6192 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2359
timestamp 1626908933
transform 1 0 6096 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1768
timestamp 1626908933
transform 1 0 6192 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_424
timestamp 1626908933
transform 1 0 6096 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3724
timestamp 1626908933
transform 1 0 6192 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1757
timestamp 1626908933
transform 1 0 6192 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3204
timestamp 1626908933
transform 1 0 6096 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1237
timestamp 1626908933
transform 1 0 6096 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3253
timestamp 1626908933
transform 1 0 6288 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1318
timestamp 1626908933
transform 1 0 6288 0 1 2553
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3203
timestamp 1626908933
transform 1 0 6096 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1236
timestamp 1626908933
transform 1 0 6096 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_593
timestamp 1626908933
transform 1 0 5760 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1315
timestamp 1626908933
transform 1 0 5760 0 1 2664
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1246
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_598
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1246
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_598
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3259
timestamp 1626908933
transform 1 0 6672 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1324
timestamp 1626908933
transform 1 0 6672 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3208
timestamp 1626908933
transform 1 0 6672 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1241
timestamp 1626908933
transform 1 0 6672 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3286
timestamp 1626908933
transform 1 0 6768 0 1 2849
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1351
timestamp 1626908933
transform 1 0 6768 0 1 2849
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_316
timestamp 1626908933
transform 1 0 7008 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_917
timestamp 1626908933
transform 1 0 7008 0 1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1265
timestamp 1626908933
transform 1 0 6864 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3232
timestamp 1626908933
transform 1 0 6864 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1349
timestamp 1626908933
transform 1 0 6864 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3284
timestamp 1626908933
transform 1 0 6864 0 1 2923
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_568
timestamp 1626908933
transform 1 0 7200 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1290
timestamp 1626908933
transform 1 0 7200 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__nand3_1  sky130_fd_sc_hs__nand3_1_0
timestamp 1626908933
transform 1 0 6528 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__nand3_1  sky130_fd_sc_hs__nand3_1_1
timestamp 1626908933
transform 1 0 6528 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_916
timestamp 1626908933
transform 1 0 7968 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_315
timestamp 1626908933
transform 1 0 7968 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1272
timestamp 1626908933
transform 1 0 8160 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_550
timestamp 1626908933
transform 1 0 8160 0 1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_859
timestamp 1626908933
transform 1 0 8592 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2794
timestamp 1626908933
transform 1 0 8592 0 1 2331
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1222
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_574
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1222
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_574
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1970
timestamp 1626908933
transform 1 0 8880 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_35
timestamp 1626908933
transform 1 0 8880 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1999
timestamp 1626908933
transform 1 0 8880 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_32
timestamp 1626908933
transform 1 0 8880 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2788
timestamp 1626908933
transform 1 0 8976 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_853
timestamp 1626908933
transform 1 0 8976 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2785
timestamp 1626908933
transform 1 0 8784 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_818
timestamp 1626908933
transform 1 0 8784 0 1 2923
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_82
timestamp 1626908933
transform 1 0 8928 0 1 2664
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_21
timestamp 1626908933
transform 1 0 8928 0 1 2664
box -38 -49 326 715
use M1M2_PR  M1M2_PR_31
timestamp 1626908933
transform 1 0 9072 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1998
timestamp 1626908933
transform 1 0 9072 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_820
timestamp 1626908933
transform 1 0 9168 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_821
timestamp 1626908933
transform 1 0 9168 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2787
timestamp 1626908933
transform 1 0 9168 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2788
timestamp 1626908933
transform 1 0 9168 0 1 2405
box -32 -32 32 32
use L1M1_PR  L1M1_PR_33
timestamp 1626908933
transform 1 0 9168 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_858
timestamp 1626908933
transform 1 0 9168 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1968
timestamp 1626908933
transform 1 0 9168 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2793
timestamp 1626908933
transform 1 0 9168 0 1 2775
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_319
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_676
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_30
timestamp 1626908933
transform 1 0 9936 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1997
timestamp 1626908933
transform 1 0 9936 0 1 2923
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_528
timestamp 1626908933
transform 1 0 9216 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1250
timestamp 1626908933
transform 1 0 9216 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_583
timestamp 1626908933
transform 1 0 10080 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1574
timestamp 1626908933
transform 1 0 10080 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2792
timestamp 1626908933
transform 1 0 10512 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_857
timestamp 1626908933
transform 1 0 10512 0 1 2405
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1573
timestamp 1626908933
transform 1 0 10560 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_582
timestamp 1626908933
transform 1 0 10560 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_825
timestamp 1626908933
transform 1 0 10704 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2792
timestamp 1626908933
transform 1 0 10704 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_863
timestamp 1626908933
transform 1 0 10704 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2798
timestamp 1626908933
transform 1 0 10704 0 1 2553
box -29 -23 29 23
use M1M2_PR  M1M2_PR_824
timestamp 1626908933
transform 1 0 10704 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2791
timestamp 1626908933
transform 1 0 10704 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_856
timestamp 1626908933
transform 1 0 10704 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2791
timestamp 1626908933
transform 1 0 10704 0 1 2775
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_680
timestamp 1626908933
transform 1 0 10656 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1671
timestamp 1626908933
transform 1 0 10656 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_427
timestamp 1626908933
transform 1 0 10176 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1025
timestamp 1626908933
transform 1 0 10176 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_15
timestamp 1626908933
transform 1 0 10752 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_77
timestamp 1626908933
transform 1 0 10752 0 1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2730
timestamp 1626908933
transform 1 0 10896 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2729
timestamp 1626908933
transform 1 0 10896 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_795
timestamp 1626908933
transform 1 0 10896 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_794
timestamp 1626908933
transform 1 0 10896 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2732
timestamp 1626908933
transform 1 0 10896 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2731
timestamp 1626908933
transform 1 0 10896 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_765
timestamp 1626908933
transform 1 0 10896 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_764
timestamp 1626908933
transform 1 0 10896 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_314
timestamp 1626908933
transform 1 0 11136 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_915
timestamp 1626908933
transform 1 0 11136 0 1 2664
box -38 -49 230 715
use L1M1_PR  L1M1_PR_862
timestamp 1626908933
transform 1 0 11088 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2797
timestamp 1626908933
transform 1 0 11088 0 1 2923
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_550
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1198
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_550
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1198
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_488
timestamp 1626908933
transform 1 0 11712 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1210
timestamp 1626908933
transform 1 0 11712 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_401
timestamp 1626908933
transform 1 0 11328 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_999
timestamp 1626908933
transform 1 0 11328 0 1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2083
timestamp 1626908933
transform 1 0 12720 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_148
timestamp 1626908933
transform 1 0 12720 0 1 2553
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2103
timestamp 1626908933
transform 1 0 12720 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2102
timestamp 1626908933
transform 1 0 12720 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_136
timestamp 1626908933
transform 1 0 12720 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_135
timestamp 1626908933
transform 1 0 12720 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_971
timestamp 1626908933
transform 1 0 12480 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_373
timestamp 1626908933
transform 1 0 12480 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_681
timestamp 1626908933
transform 1 0 12864 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1672
timestamp 1626908933
transform 1 0 12864 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_147
timestamp 1626908933
transform 1 0 13008 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2082
timestamp 1626908933
transform 1 0 13008 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_581
timestamp 1626908933
transform 1 0 13536 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1572
timestamp 1626908933
transform 1 0 13536 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_973
timestamp 1626908933
transform 1 0 13296 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1608
timestamp 1626908933
transform 1 0 13488 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2908
timestamp 1626908933
transform 1 0 13296 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3543
timestamp 1626908933
transform 1 0 13488 0 1 2775
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_14
timestamp 1626908933
transform -1 0 13536 0 1 2664
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_53
timestamp 1626908933
transform -1 0 13536 0 1 2664
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1174
timestamp 1626908933
transform 1 0 13700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_526
timestamp 1626908933
transform 1 0 13700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1174
timestamp 1626908933
transform 1 0 13700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_526
timestamp 1626908933
transform 1 0 13700 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1171
timestamp 1626908933
transform 1 0 13632 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_449
timestamp 1626908933
transform 1 0 13632 0 1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_920
timestamp 1626908933
transform 1 0 13872 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2887
timestamp 1626908933
transform 1 0 13872 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_313
timestamp 1626908933
transform 1 0 14400 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_914
timestamp 1626908933
transform 1 0 14400 0 1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1714
timestamp 1626908933
transform 1 0 14352 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1938
timestamp 1626908933
transform 1 0 14544 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3681
timestamp 1626908933
transform 1 0 14352 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3905
timestamp 1626908933
transform 1 0 14544 0 1 2405
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1904
timestamp 1626908933
transform 1 0 14544 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3839
timestamp 1626908933
transform 1 0 14544 0 1 2405
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_337
timestamp 1626908933
transform 1 0 14592 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_935
timestamp 1626908933
transform 1 0 14592 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_318
timestamp 1626908933
transform 1 0 14976 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_675
timestamp 1626908933
transform 1 0 14976 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1520
timestamp 1626908933
transform 1 0 14736 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1521
timestamp 1626908933
transform 1 0 14736 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3487
timestamp 1626908933
transform 1 0 14736 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3488
timestamp 1626908933
transform 1 0 14736 0 1 2405
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1607
timestamp 1626908933
transform 1 0 14832 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3542
timestamp 1626908933
transform 1 0 14832 0 1 2405
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_580
timestamp 1626908933
transform 1 0 15456 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1571
timestamp 1626908933
transform 1 0 15456 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_47
timestamp 1626908933
transform 1 0 15216 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1982
timestamp 1626908933
transform 1 0 15216 0 1 2553
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_324
timestamp 1626908933
transform 1 0 15072 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_922
timestamp 1626908933
transform 1 0 15072 0 1 2664
box -38 -49 422 715
use M1M2_PR  M1M2_PR_42
timestamp 1626908933
transform 1 0 15792 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_43
timestamp 1626908933
transform 1 0 15792 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2009
timestamp 1626908933
transform 1 0 15792 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2010
timestamp 1626908933
transform 1 0 15792 0 1 2553
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_579
timestamp 1626908933
transform 1 0 16320 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1570
timestamp 1626908933
transform 1 0 16320 0 1 2664
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_502
timestamp 1626908933
transform 1 0 16100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1150
timestamp 1626908933
transform 1 0 16100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_502
timestamp 1626908933
transform 1 0 16100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1150
timestamp 1626908933
transform 1 0 16100 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_416
timestamp 1626908933
transform 1 0 15552 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1138
timestamp 1626908933
transform 1 0 15552 0 1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1980
timestamp 1626908933
transform 1 0 16464 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_45
timestamp 1626908933
transform 1 0 16464 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_19
timestamp 1626908933
transform 1 0 16416 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_88
timestamp 1626908933
transform 1 0 16416 0 1 2664
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3836
timestamp 1626908933
transform 1 0 17040 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1901
timestamp 1626908933
transform 1 0 17040 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1569
timestamp 1626908933
transform 1 0 16896 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_578
timestamp 1626908933
transform 1 0 16896 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1092
timestamp 1626908933
transform 1 0 16992 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_370
timestamp 1626908933
transform 1 0 16992 0 1 2664
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1126
timestamp 1626908933
transform 1 0 18500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_478
timestamp 1626908933
transform 1 0 18500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1126
timestamp 1626908933
transform 1 0 18500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_478
timestamp 1626908933
transform 1 0 18500 0 1 2664
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3835
timestamp 1626908933
transform 1 0 18096 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1900
timestamp 1626908933
transform 1 0 18096 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3901
timestamp 1626908933
transform 1 0 18096 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1934
timestamp 1626908933
transform 1 0 18096 0 1 2923
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_48
timestamp 1626908933
transform 1 0 17760 0 1 2664
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_23
timestamp 1626908933
transform 1 0 17760 0 1 2664
box -38 -49 2246 715
use M1M2_PR  M1M2_PR_3663
timestamp 1626908933
transform 1 0 19440 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3661
timestamp 1626908933
transform 1 0 19536 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1696
timestamp 1626908933
transform 1 0 19440 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1694
timestamp 1626908933
transform 1 0 19536 0 1 2331
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1033
timestamp 1626908933
transform 1 0 20064 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_311
timestamp 1626908933
transform 1 0 20064 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_674
timestamp 1626908933
transform 1 0 19968 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_317
timestamp 1626908933
transform 1 0 19968 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1928
timestamp 1626908933
transform 1 0 20400 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1929
timestamp 1626908933
transform 1 0 20400 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3895
timestamp 1626908933
transform 1 0 20400 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3896
timestamp 1626908933
transform 1 0 20400 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1897
timestamp 1626908933
transform 1 0 20400 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3832
timestamp 1626908933
transform 1 0 20400 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_372
timestamp 1626908933
transform 1 0 20832 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_973
timestamp 1626908933
transform 1 0 20832 0 1 2664
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_454
timestamp 1626908933
transform 1 0 20900 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1102
timestamp 1626908933
transform 1 0 20900 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_454
timestamp 1626908933
transform 1 0 20900 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1102
timestamp 1626908933
transform 1 0 20900 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_96
timestamp 1626908933
transform 1 0 21024 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_27
timestamp 1626908933
transform 1 0 21024 0 1 2664
box -38 -49 518 715
use M1M2_PR  M1M2_PR_105
timestamp 1626908933
transform 1 0 21168 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_106
timestamp 1626908933
transform 1 0 21168 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_796
timestamp 1626908933
transform 1 0 21456 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2072
timestamp 1626908933
transform 1 0 21168 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2073
timestamp 1626908933
transform 1 0 21168 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2763
timestamp 1626908933
transform 1 0 21456 0 1 2997
box -32 -32 32 32
use L1M1_PR  L1M1_PR_119
timestamp 1626908933
transform 1 0 21168 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2054
timestamp 1626908933
transform 1 0 21168 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_577
timestamp 1626908933
transform 1 0 21504 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1568
timestamp 1626908933
transform 1 0 21504 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_193
timestamp 1626908933
transform 1 0 21600 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_791
timestamp 1626908933
transform 1 0 21600 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_997
timestamp 1626908933
transform 1 0 21984 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_275
timestamp 1626908933
transform 1 0 21984 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_98
timestamp 1626908933
transform -1 0 23136 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_36
timestamp 1626908933
transform -1 0 23136 0 1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2052
timestamp 1626908933
transform 1 0 22224 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_117
timestamp 1626908933
transform 1 0 22224 0 1 2553
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_576
timestamp 1626908933
transform 1 0 23136 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1567
timestamp 1626908933
transform 1 0 23136 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_827
timestamp 1626908933
transform 1 0 22992 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2762
timestamp 1626908933
transform 1 0 22992 0 1 2997
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_430
timestamp 1626908933
transform 1 0 23300 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1078
timestamp 1626908933
transform 1 0 23300 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_430
timestamp 1626908933
transform 1 0 23300 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1078
timestamp 1626908933
transform 1 0 23300 0 1 2664
box -100 -49 100 49
use M1M2_PR  M1M2_PR_101
timestamp 1626908933
transform 1 0 23664 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2068
timestamp 1626908933
transform 1 0 23664 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_236
timestamp 1626908933
transform 1 0 23232 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_958
timestamp 1626908933
transform 1 0 23232 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_312
timestamp 1626908933
transform 1 0 24000 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_913
timestamp 1626908933
transform 1 0 24000 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_575
timestamp 1626908933
transform 1 0 24192 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1566
timestamp 1626908933
transform 1 0 24192 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_113
timestamp 1626908933
transform 1 0 24336 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2048
timestamp 1626908933
transform 1 0 24336 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_3
timestamp 1626908933
transform 1 0 24288 0 1 2664
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_65
timestamp 1626908933
transform 1 0 24288 0 1 2664
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_10
timestamp 1626908933
transform 1 0 24576 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_62
timestamp 1626908933
transform 1 0 24576 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_316
timestamp 1626908933
transform 1 0 24960 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_673
timestamp 1626908933
transform 1 0 24960 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_574
timestamp 1626908933
transform 1 0 25056 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1565
timestamp 1626908933
transform 1 0 25056 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_112
timestamp 1626908933
transform 1 0 26112 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_710
timestamp 1626908933
transform 1 0 26112 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_311
timestamp 1626908933
transform 1 0 25920 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_912
timestamp 1626908933
transform 1 0 25920 0 1 2664
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_406
timestamp 1626908933
transform 1 0 25700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1054
timestamp 1626908933
transform 1 0 25700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_406
timestamp 1626908933
transform 1 0 25700 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1054
timestamp 1626908933
transform 1 0 25700 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_195
timestamp 1626908933
transform 1 0 25152 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_917
timestamp 1626908933
transform 1 0 25152 0 1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1923
timestamp 1626908933
transform 1 0 26832 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1924
timestamp 1626908933
transform 1 0 26832 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3890
timestamp 1626908933
transform 1 0 26832 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3891
timestamp 1626908933
transform 1 0 26832 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1892
timestamp 1626908933
transform 1 0 26832 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3827
timestamp 1626908933
transform 1 0 26832 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_573
timestamp 1626908933
transform 1 0 27264 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_682
timestamp 1626908933
transform 1 0 27360 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1564
timestamp 1626908933
transform 1 0 27264 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1673
timestamp 1626908933
transform 1 0 27360 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1684
timestamp 1626908933
transform 1 0 27024 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1776
timestamp 1626908933
transform 1 0 27120 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3651
timestamp 1626908933
transform 1 0 27024 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3743
timestamp 1626908933
transform 1 0 27120 0 1 2553
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_167
timestamp 1626908933
transform 1 0 26496 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_889
timestamp 1626908933
transform 1 0 26496 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_46
timestamp 1626908933
transform 1 0 27456 0 1 2664
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_21
timestamp 1626908933
transform 1 0 27456 0 1 2664
box -38 -49 2246 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_382
timestamp 1626908933
transform 1 0 28100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1030
timestamp 1626908933
transform 1 0 28100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_382
timestamp 1626908933
transform 1 0 28100 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1030
timestamp 1626908933
transform 1 0 28100 0 1 2664
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1683
timestamp 1626908933
transform 1 0 27696 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1922
timestamp 1626908933
transform 1 0 27888 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3650
timestamp 1626908933
transform 1 0 27696 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3889
timestamp 1626908933
transform 1 0 27888 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1891
timestamp 1626908933
transform 1 0 27792 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3826
timestamp 1626908933
transform 1 0 27792 0 1 2923
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1674
timestamp 1626908933
transform 1 0 29856 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_683
timestamp 1626908933
transform 1 0 29856 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_974
timestamp 1626908933
transform 1 0 29664 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_911
timestamp 1626908933
transform 1 0 30048 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_373
timestamp 1626908933
transform 1 0 29664 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_310
timestamp 1626908933
transform 1 0 30048 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_672
timestamp 1626908933
transform 1 0 29952 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_315
timestamp 1626908933
transform 1 0 29952 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3746
timestamp 1626908933
transform 1 0 30288 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1779
timestamp 1626908933
transform 1 0 30288 0 1 2923
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1563
timestamp 1626908933
transform 1 0 30240 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_572
timestamp 1626908933
transform 1 0 30240 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_786
timestamp 1626908933
transform 1 0 30336 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_64
timestamp 1626908933
transform 1 0 30336 0 1 2664
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1006
timestamp 1626908933
transform 1 0 30500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_358
timestamp 1626908933
transform 1 0 30500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1006
timestamp 1626908933
transform 1 0 30500 0 1 2664
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_358
timestamp 1626908933
transform 1 0 30500 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1562
timestamp 1626908933
transform 1 0 31104 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_571
timestamp 1626908933
transform 1 0 31104 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_743
timestamp 1626908933
transform 1 0 31200 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_21
timestamp 1626908933
transform 1 0 31200 0 1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3744
timestamp 1626908933
transform 1 0 31920 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3741
timestamp 1626908933
transform 1 0 32016 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1777
timestamp 1626908933
transform 1 0 31920 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1774
timestamp 1626908933
transform 1 0 32016 0 1 2553
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1675
timestamp 1626908933
transform 1 0 31968 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_684
timestamp 1626908933
transform 1 0 31968 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_309
timestamp 1626908933
transform 1 0 0 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_910
timestamp 1626908933
transform 1 0 0 0 -1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1958
timestamp 1626908933
transform 1 0 144 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3925
timestamp 1626908933
transform 1 0 144 0 1 3515
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_333
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_981
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_333
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_981
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_719
timestamp 1626908933
transform 1 0 192 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1441
timestamp 1626908933
transform 1 0 192 0 -1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3212
timestamp 1626908933
transform 1 0 1584 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1245
timestamp 1626908933
transform 1 0 1584 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1561
timestamp 1626908933
transform 1 0 960 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_570
timestamp 1626908933
transform 1 0 960 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1180
timestamp 1626908933
transform 1 0 1056 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_582
timestamp 1626908933
transform 1 0 1056 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1408
timestamp 1626908933
transform 1 0 1440 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_686
timestamp 1626908933
transform 1 0 1440 0 -1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3224
timestamp 1626908933
transform 1 0 2448 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1257
timestamp 1626908933
transform 1 0 2448 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1560
timestamp 1626908933
transform 1 0 2208 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_569
timestamp 1626908933
transform 1 0 2208 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_975
timestamp 1626908933
transform 1 0 2304 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_374
timestamp 1626908933
transform 1 0 2304 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_671
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_314
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_10
timestamp 1626908933
transform 1 0 2688 0 -1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_4
timestamp 1626908933
transform 1 0 2688 0 -1 3996
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3263
timestamp 1626908933
transform 1 0 2736 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1328
timestamp 1626908933
transform 1 0 2736 0 1 3737
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1676
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_685
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_957
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_309
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_957
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_309
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3275
timestamp 1626908933
transform 1 0 2928 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3257
timestamp 1626908933
transform 1 0 3024 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1340
timestamp 1626908933
transform 1 0 2928 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1322
timestamp 1626908933
transform 1 0 3024 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3207
timestamp 1626908933
transform 1 0 2832 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1240
timestamp 1626908933
transform 1 0 2832 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_909
timestamp 1626908933
transform 1 0 3168 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_308
timestamp 1626908933
transform 1 0 3168 0 -1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1235
timestamp 1626908933
transform 1 0 3312 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3202
timestamp 1626908933
transform 1 0 3312 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_649
timestamp 1626908933
transform 1 0 3360 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1371
timestamp 1626908933
transform 1 0 3360 0 -1 3996
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3251
timestamp 1626908933
transform 1 0 4272 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1316
timestamp 1626908933
transform 1 0 4272 0 1 3219
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_976
timestamp 1626908933
transform 1 0 4320 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_908
timestamp 1626908933
transform 1 0 4128 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_375
timestamp 1626908933
transform 1 0 4320 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_307
timestamp 1626908933
transform 1 0 4128 0 -1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3862
timestamp 1626908933
transform 1 0 4464 0 1 3515
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3241
timestamp 1626908933
transform 1 0 4752 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1927
timestamp 1626908933
transform 1 0 4464 0 1 3515
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1306
timestamp 1626908933
transform 1 0 4752 0 1 3737
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3922
timestamp 1626908933
transform 1 0 4560 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3196
timestamp 1626908933
transform 1 0 4656 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1955
timestamp 1626908933
transform 1 0 4560 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1229
timestamp 1626908933
transform 1 0 4656 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_907
timestamp 1626908933
transform 1 0 4800 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_306
timestamp 1626908933
transform 1 0 4800 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_115
timestamp 1626908933
transform 1 0 4512 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_54
timestamp 1626908933
transform 1 0 4512 0 -1 3996
box -38 -49 326 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_285
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_933
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_285
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_933
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_611
timestamp 1626908933
transform 1 0 4992 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1333
timestamp 1626908933
transform 1 0 4992 0 -1 3996
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3255
timestamp 1626908933
transform 1 0 5328 0 1 3145
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1320
timestamp 1626908933
transform 1 0 5328 0 1 3145
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3285
timestamp 1626908933
transform 1 0 6096 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3240
timestamp 1626908933
transform 1 0 5904 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2284
timestamp 1626908933
transform 1 0 6096 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1350
timestamp 1626908933
transform 1 0 6096 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1305
timestamp 1626908933
transform 1 0 5904 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_349
timestamp 1626908933
transform 1 0 6096 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2290
timestamp 1626908933
transform 1 0 6192 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_323
timestamp 1626908933
transform 1 0 6192 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_6
timestamp 1626908933
transform -1 0 6240 0 -1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_14
timestamp 1626908933
transform -1 0 6240 0 -1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1559
timestamp 1626908933
transform 1 0 6432 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_568
timestamp 1626908933
transform 1 0 6432 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_906
timestamp 1626908933
transform 1 0 6240 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_305
timestamp 1626908933
transform 1 0 6240 0 -1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3232
timestamp 1626908933
transform 1 0 6672 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1297
timestamp 1626908933
transform 1 0 6672 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3190
timestamp 1626908933
transform 1 0 6672 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1223
timestamp 1626908933
transform 1 0 6672 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3231
timestamp 1626908933
transform 1 0 6864 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1264
timestamp 1626908933
transform 1 0 6864 0 1 3441
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_582
timestamp 1626908933
transform 1 0 6528 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1304
timestamp 1626908933
transform 1 0 6528 0 -1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1525
timestamp 1626908933
transform 1 0 6960 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3492
timestamp 1626908933
transform 1 0 6960 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_567
timestamp 1626908933
transform 1 0 7296 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1558
timestamp 1626908933
transform 1 0 7296 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_313
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_670
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_686
timestamp 1626908933
transform 1 0 7392 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1677
timestamp 1626908933
transform 1 0 7392 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1611
timestamp 1626908933
transform 1 0 7632 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3546
timestamp 1626908933
transform 1 0 7632 0 1 3737
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_261
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_909
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_261
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_909
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1748
timestamp 1626908933
transform 1 0 7824 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3715
timestamp 1626908933
transform 1 0 7824 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1942
timestamp 1626908933
transform 1 0 7920 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3909
timestamp 1626908933
transform 1 0 7920 0 1 3737
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1912
timestamp 1626908933
transform 1 0 7920 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3847
timestamp 1626908933
transform 1 0 7920 0 1 3737
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_28
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_3
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1249
timestamp 1626908933
transform 1 0 9792 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_527
timestamp 1626908933
transform 1 0 9792 0 -1 3996
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_885
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_237
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_885
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_237
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3694
timestamp 1626908933
transform 1 0 10320 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1727
timestamp 1626908933
transform 1 0 10320 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1007
timestamp 1626908933
transform 1 0 10560 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_409
timestamp 1626908933
transform 1 0 10560 0 -1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3440
timestamp 1626908933
transform 1 0 10992 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1473
timestamp 1626908933
transform 1 0 10992 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1557
timestamp 1626908933
transform 1 0 10944 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_566
timestamp 1626908933
transform 1 0 10944 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1220
timestamp 1626908933
transform 1 0 11040 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_498
timestamp 1626908933
transform 1 0 11040 0 -1 3996
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3494
timestamp 1626908933
transform 1 0 11088 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1559
timestamp 1626908933
transform 1 0 11088 0 1 3219
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_905
timestamp 1626908933
transform 1 0 11808 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_304
timestamp 1626908933
transform 1 0 11808 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_565
timestamp 1626908933
transform 1 0 12000 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1556
timestamp 1626908933
transform 1 0 12000 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_312
timestamp 1626908933
transform 1 0 12480 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_669
timestamp 1626908933
transform 1 0 12480 0 -1 3996
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_213
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_861
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_213
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_861
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_366
timestamp 1626908933
transform 1 0 12576 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_382
timestamp 1626908933
transform 1 0 12096 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_964
timestamp 1626908933
transform 1 0 12576 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_980
timestamp 1626908933
transform 1 0 12096 0 -1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2902
timestamp 1626908933
transform 1 0 13104 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_967
timestamp 1626908933
transform 1 0 13104 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2881
timestamp 1626908933
transform 1 0 13104 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_914
timestamp 1626908933
transform 1 0 13104 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1187
timestamp 1626908933
transform 1 0 12960 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_465
timestamp 1626908933
transform 1 0 12960 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_904
timestamp 1626908933
transform 1 0 13728 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_303
timestamp 1626908933
transform 1 0 13728 0 -1 3996
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_189
timestamp 1626908933
transform 1 0 14900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_837
timestamp 1626908933
transform 1 0 14900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_189
timestamp 1626908933
transform 1 0 14900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_837
timestamp 1626908933
transform 1 0 14900 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1519
timestamp 1626908933
transform 1 0 14832 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1713
timestamp 1626908933
transform 1 0 14352 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3486
timestamp 1626908933
transform 1 0 14832 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3680
timestamp 1626908933
transform 1 0 14352 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1605
timestamp 1626908933
transform 1 0 14736 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1903
timestamp 1626908933
transform 1 0 15024 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3540
timestamp 1626908933
transform 1 0 14736 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3838
timestamp 1626908933
transform 1 0 15024 0 1 3737
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_434
timestamp 1626908933
transform 1 0 13920 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1156
timestamp 1626908933
transform 1 0 13920 0 -1 3996
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2676
timestamp 1626908933
transform 1 0 16560 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_741
timestamp 1626908933
transform 1 0 16560 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2684
timestamp 1626908933
transform 1 0 16464 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_717
timestamp 1626908933
transform 1 0 16464 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_31
timestamp 1626908933
transform 1 0 14688 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_6
timestamp 1626908933
transform 1 0 14688 0 -1 3996
box -38 -49 2246 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_813
timestamp 1626908933
transform 1 0 17300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_165
timestamp 1626908933
transform 1 0 17300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_813
timestamp 1626908933
transform 1 0 17300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_165
timestamp 1626908933
transform 1 0 17300 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_977
timestamp 1626908933
transform 1 0 17280 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_376
timestamp 1626908933
transform 1 0 17280 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_887
timestamp 1626908933
transform 1 0 16896 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_289
timestamp 1626908933
transform 1 0 16896 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_311
timestamp 1626908933
transform 1 0 17472 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_668
timestamp 1626908933
transform 1 0 17472 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1572
timestamp 1626908933
transform 1 0 17808 0 1 3071
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3507
timestamp 1626908933
transform 1 0 17808 0 1 3071
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1484
timestamp 1626908933
transform 1 0 17904 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1485
timestamp 1626908933
transform 1 0 17904 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3451
timestamp 1626908933
transform 1 0 17904 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3452
timestamp 1626908933
transform 1 0 17904 0 1 3071
box -32 -32 32 32
use L1M1_PR  L1M1_PR_946
timestamp 1626908933
transform 1 0 18192 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1571
timestamp 1626908933
transform 1 0 18000 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2881
timestamp 1626908933
transform 1 0 18192 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3506
timestamp 1626908933
transform 1 0 18000 0 1 3441
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_274
timestamp 1626908933
transform 1 0 17568 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_872
timestamp 1626908933
transform 1 0 17568 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_23
timestamp 1626908933
transform 1 0 17952 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_62
timestamp 1626908933
transform 1 0 17952 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_302
timestamp 1626908933
transform 1 0 18528 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_903
timestamp 1626908933
transform 1 0 18528 0 -1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_190
timestamp 1626908933
transform 1 0 18672 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_898
timestamp 1626908933
transform 1 0 18288 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2157
timestamp 1626908933
transform 1 0 18672 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2865
timestamp 1626908933
transform 1 0 18288 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1040
timestamp 1626908933
transform 1 0 18384 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2975
timestamp 1626908933
transform 1 0 18384 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_977
timestamp 1626908933
transform 1 0 18864 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2944
timestamp 1626908933
transform 1 0 18864 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_340
timestamp 1626908933
transform 1 0 18720 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1062
timestamp 1626908933
transform 1 0 18720 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_301
timestamp 1626908933
transform 1 0 19488 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_902
timestamp 1626908933
transform 1 0 19488 0 -1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1695
timestamp 1626908933
transform 1 0 19440 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3662
timestamp 1626908933
transform 1 0 19440 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_687
timestamp 1626908933
transform 1 0 19680 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1678
timestamp 1626908933
transform 1 0 19680 0 -1 3996
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_141
timestamp 1626908933
transform 1 0 19700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_789
timestamp 1626908933
transform 1 0 19700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_141
timestamp 1626908933
transform 1 0 19700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_789
timestamp 1626908933
transform 1 0 19700 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_206
timestamp 1626908933
transform 1 0 19920 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2141
timestamp 1626908933
transform 1 0 19920 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1927
timestamp 1626908933
transform 1 0 20400 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3894
timestamp 1626908933
transform 1 0 20400 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_738
timestamp 1626908933
transform 1 0 20976 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2705
timestamp 1626908933
transform 1 0 20976 0 1 3219
box -32 -32 32 32
use L1M1_PR  L1M1_PR_759
timestamp 1626908933
transform 1 0 21168 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2694
timestamp 1626908933
transform 1 0 21168 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1896
timestamp 1626908933
transform 1 0 21648 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3831
timestamp 1626908933
transform 1 0 21648 0 1 3737
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_765
timestamp 1626908933
transform 1 0 22100 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_117
timestamp 1626908933
transform 1 0 22100 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_765
timestamp 1626908933
transform 1 0 22100 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_117
timestamp 1626908933
transform 1 0 22100 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3509
timestamp 1626908933
transform 1 0 21936 0 1 3589
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1574
timestamp 1626908933
transform 1 0 21936 0 1 3589
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1555
timestamp 1626908933
transform 1 0 21984 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_564
timestamp 1626908933
transform 1 0 21984 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_786
timestamp 1626908933
transform 1 0 22080 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_188
timestamp 1626908933
transform 1 0 22080 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_47
timestamp 1626908933
transform -1 0 21984 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_22
timestamp 1626908933
transform -1 0 21984 0 -1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_310
timestamp 1626908933
transform 1 0 22464 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_667
timestamp 1626908933
transform 1 0 22464 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3508
timestamp 1626908933
transform 1 0 22800 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2973
timestamp 1626908933
transform 1 0 22704 0 1 3145
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1573
timestamp 1626908933
transform 1 0 22800 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1038
timestamp 1626908933
transform 1 0 22704 0 1 3145
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3454
timestamp 1626908933
transform 1 0 22800 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2942
timestamp 1626908933
transform 1 0 22704 0 1 3145
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1487
timestamp 1626908933
transform 1 0 22800 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_975
timestamp 1626908933
transform 1 0 22704 0 1 3145
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3453
timestamp 1626908933
transform 1 0 22800 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2941
timestamp 1626908933
transform 1 0 22704 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1486
timestamp 1626908933
transform 1 0 22800 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_974
timestamp 1626908933
transform 1 0 22704 0 1 3441
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_90
timestamp 1626908933
transform 1 0 22944 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_28
timestamp 1626908933
transform 1 0 22944 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_11
timestamp 1626908933
transform 1 0 22560 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_63
timestamp 1626908933
transform 1 0 22560 0 -1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_578
timestamp 1626908933
transform 1 0 22992 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_973
timestamp 1626908933
transform 1 0 23184 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2545
timestamp 1626908933
transform 1 0 22992 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2940
timestamp 1626908933
transform 1 0 23184 0 1 3219
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1036
timestamp 1626908933
transform 1 0 23184 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2971
timestamp 1626908933
transform 1 0 23184 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_972
timestamp 1626908933
transform 1 0 23184 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2939
timestamp 1626908933
transform 1 0 23184 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1035
timestamp 1626908933
transform 1 0 23184 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1037
timestamp 1626908933
transform 1 0 23088 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2970
timestamp 1626908933
transform 1 0 23184 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2972
timestamp 1626908933
transform 1 0 23088 0 1 3441
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_235
timestamp 1626908933
transform 1 0 23232 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_957
timestamp 1626908933
transform 1 0 23232 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1554
timestamp 1626908933
transform 1 0 24384 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_563
timestamp 1626908933
transform 1 0 24384 0 -1 3996
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_741
timestamp 1626908933
transform 1 0 24500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_93
timestamp 1626908933
transform 1 0 24500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_741
timestamp 1626908933
transform 1 0 24500 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_93
timestamp 1626908933
transform 1 0 24500 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2681
timestamp 1626908933
transform 1 0 24624 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2516
timestamp 1626908933
transform 1 0 24432 0 1 3145
box -29 -23 29 23
use L1M1_PR  L1M1_PR_746
timestamp 1626908933
transform 1 0 24624 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_581
timestamp 1626908933
transform 1 0 24432 0 1 3145
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_205
timestamp 1626908933
transform 1 0 24480 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_927
timestamp 1626908933
transform 1 0 24480 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_146
timestamp 1626908933
transform 1 0 24000 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_744
timestamp 1626908933
transform 1 0 24000 0 -1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2688
timestamp 1626908933
transform 1 0 24720 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_721
timestamp 1626908933
transform 1 0 24720 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_717
timestamp 1626908933
transform 1 0 25248 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_119
timestamp 1626908933
transform 1 0 25248 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_10
timestamp 1626908933
transform -1 0 26112 0 -1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_79
timestamp 1626908933
transform -1 0 26112 0 -1 3996
box -38 -49 518 715
use M1M2_PR  M1M2_PR_2938
timestamp 1626908933
transform 1 0 25968 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_971
timestamp 1626908933
transform 1 0 25968 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_59
timestamp 1626908933
transform 1 0 26112 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_7
timestamp 1626908933
transform 1 0 26112 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_888
timestamp 1626908933
transform 1 0 26496 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_166
timestamp 1626908933
transform 1 0 26496 0 -1 3996
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_717
timestamp 1626908933
transform 1 0 26900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_69
timestamp 1626908933
transform 1 0 26900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_717
timestamp 1626908933
transform 1 0 26900 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_69
timestamp 1626908933
transform 1 0 26900 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_978
timestamp 1626908933
transform 1 0 27264 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_377
timestamp 1626908933
transform 1 0 27264 0 -1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3511
timestamp 1626908933
transform 1 0 27504 0 1 3071
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1576
timestamp 1626908933
transform 1 0 27504 0 1 3071
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_901
timestamp 1626908933
transform 1 0 27552 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_300
timestamp 1626908933
transform 1 0 27552 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_666
timestamp 1626908933
transform 1 0 27456 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_309
timestamp 1626908933
transform 1 0 27456 0 -1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3456
timestamp 1626908933
transform 1 0 28272 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1489
timestamp 1626908933
transform 1 0 28272 0 1 3071
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_857
timestamp 1626908933
transform 1 0 27744 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_135
timestamp 1626908933
transform 1 0 27744 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_562
timestamp 1626908933
transform 1 0 28896 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1553
timestamp 1626908933
transform 1 0 28896 0 -1 3996
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_45
timestamp 1626908933
transform 1 0 29300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_693
timestamp 1626908933
transform 1 0 29300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_45
timestamp 1626908933
transform 1 0 29300 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_693
timestamp 1626908933
transform 1 0 29300 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_100
timestamp 1626908933
transform 1 0 28992 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_822
timestamp 1626908933
transform 1 0 28992 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_67
timestamp 1626908933
transform 1 0 28512 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_665
timestamp 1626908933
transform 1 0 28512 0 -1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2134
timestamp 1626908933
transform 1 0 29616 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_199
timestamp 1626908933
transform 1 0 29616 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2150
timestamp 1626908933
transform 1 0 29616 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_183
timestamp 1626908933
transform 1 0 29616 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_900
timestamp 1626908933
transform 1 0 29760 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_299
timestamp 1626908933
transform 1 0 29760 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_634
timestamp 1626908933
transform 1 0 29952 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_36
timestamp 1626908933
transform 1 0 29952 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_785
timestamp 1626908933
transform 1 0 30336 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_63
timestamp 1626908933
transform 1 0 30336 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_612
timestamp 1626908933
transform 1 0 31104 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_14
timestamp 1626908933
transform 1 0 31104 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_561
timestamp 1626908933
transform 1 0 31488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1552
timestamp 1626908933
transform 1 0 31488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_308
timestamp 1626908933
transform 1 0 31680 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_665
timestamp 1626908933
transform 1 0 31680 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_688
timestamp 1626908933
transform 1 0 31584 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1679
timestamp 1626908933
transform 1 0 31584 0 -1 3996
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_21
timestamp 1626908933
transform 1 0 31700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_669
timestamp 1626908933
transform 1 0 31700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_21
timestamp 1626908933
transform 1 0 31700 0 1 3330
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_669
timestamp 1626908933
transform 1 0 31700 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_378
timestamp 1626908933
transform 1 0 31776 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_979
timestamp 1626908933
transform 1 0 31776 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1680
timestamp 1626908933
transform 1 0 31968 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_689
timestamp 1626908933
transform 1 0 31968 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_307
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_664
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_379
timestamp 1626908933
transform 1 0 0 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_980
timestamp 1626908933
transform 1 0 0 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_690
timestamp 1626908933
transform 1 0 192 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1681
timestamp 1626908933
transform 1 0 192 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1954
timestamp 1626908933
transform 1 0 144 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3921
timestamp 1626908933
transform 1 0 144 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_691
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1682
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1923
timestamp 1626908933
transform 1 0 528 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3858
timestamp 1626908933
transform 1 0 528 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_135
timestamp 1626908933
transform 1 0 480 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_66
timestamp 1626908933
transform 1 0 480 0 1 3996
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1342
timestamp 1626908933
transform 1 0 1008 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3277
timestamp 1626908933
transform 1 0 1008 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1247
timestamp 1626908933
transform 1 0 1488 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3214
timestamp 1626908933
transform 1 0 1488 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1327
timestamp 1626908933
transform 1 0 1488 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3262
timestamp 1626908933
transform 1 0 1488 0 1 4551
box -29 -23 29 23
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_3
timestamp 1626908933
transform -1 0 1632 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_8
timestamp 1626908933
transform -1 0 1632 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_12
timestamp 1626908933
transform 1 0 960 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_64
timestamp 1626908933
transform 1 0 960 0 1 3996
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1293
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_645
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1293
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_645
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3265
timestamp 1626908933
transform 1 0 1776 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1330
timestamp 1626908933
transform 1 0 1776 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1683
timestamp 1626908933
transform 1 0 1824 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_692
timestamp 1626908933
transform 1 0 1824 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_981
timestamp 1626908933
transform 1 0 1632 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_380
timestamp 1626908933
transform 1 0 1632 0 1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1243
timestamp 1626908933
transform 1 0 1872 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3210
timestamp 1626908933
transform 1 0 1872 0 1 4551
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1329
timestamp 1626908933
transform 1 0 2064 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1341
timestamp 1626908933
transform 1 0 2160 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3264
timestamp 1626908933
transform 1 0 2064 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3276
timestamp 1626908933
transform 1 0 2160 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_13
timestamp 1626908933
transform -1 0 2400 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_5
timestamp 1626908933
transform -1 0 2400 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_381
timestamp 1626908933
transform 1 0 2400 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_982
timestamp 1626908933
transform 1 0 2400 0 1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1256
timestamp 1626908933
transform 1 0 2448 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3223
timestamp 1626908933
transform 1 0 2448 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1323
timestamp 1626908933
transform 1 0 2256 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3258
timestamp 1626908933
transform 1 0 2256 0 1 4403
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1253
timestamp 1626908933
transform 1 0 2736 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3220
timestamp 1626908933
transform 1 0 2736 0 1 4551
box -32 -32 32 32
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_5
timestamp 1626908933
transform -1 0 3264 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_13
timestamp 1626908933
transform -1 0 3264 0 1 3996
box -38 -49 710 715
use M1M2_PR  M1M2_PR_1255
timestamp 1626908933
transform 1 0 3024 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3222
timestamp 1626908933
transform 1 0 3024 0 1 3885
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1338
timestamp 1626908933
transform 1 0 3120 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3273
timestamp 1626908933
transform 1 0 3120 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3274
timestamp 1626908933
transform 1 0 2928 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1339
timestamp 1626908933
transform 1 0 2928 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3221
timestamp 1626908933
transform 1 0 3024 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1254
timestamp 1626908933
transform 1 0 3024 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3233
timestamp 1626908933
transform 1 0 3504 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1266
timestamp 1626908933
transform 1 0 3504 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3206
timestamp 1626908933
transform 1 0 2832 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1239
timestamp 1626908933
transform 1 0 2832 0 1 4403
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2281
timestamp 1626908933
transform 1 0 2928 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_346
timestamp 1626908933
transform 1 0 2928 0 1 4403
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2287
timestamp 1626908933
transform 1 0 3120 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_320
timestamp 1626908933
transform 1 0 3120 0 1 4403
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3272
timestamp 1626908933
transform 1 0 2832 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1337
timestamp 1626908933
transform 1 0 2832 0 1 4551
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_540
timestamp 1626908933
transform 1 0 3264 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1138
timestamp 1626908933
transform 1 0 3264 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_560
timestamp 1626908933
transform 1 0 3936 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1551
timestamp 1626908933
transform 1 0 3936 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1307
timestamp 1626908933
transform 1 0 3792 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1354
timestamp 1626908933
transform 1 0 3696 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3242
timestamp 1626908933
transform 1 0 3792 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3289
timestamp 1626908933
transform 1 0 3696 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_2
timestamp 1626908933
transform 1 0 3648 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_7
timestamp 1626908933
transform 1 0 3648 0 1 3996
box -38 -49 326 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_621
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1269
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_621
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1269
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_632
timestamp 1626908933
transform 1 0 4032 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1354
timestamp 1626908933
transform 1 0 4032 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_559
timestamp 1626908933
transform 1 0 4800 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1550
timestamp 1626908933
transform 1 0 4800 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1228
timestamp 1626908933
transform 1 0 4656 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3195
timestamp 1626908933
transform 1 0 4656 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1304
timestamp 1626908933
transform 1 0 4752 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3239
timestamp 1626908933
transform 1 0 4752 0 1 3885
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_306
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_663
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_298
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_899
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_693
timestamp 1626908933
transform 1 0 4896 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1684
timestamp 1626908933
transform 1 0 4896 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1227
timestamp 1626908933
transform 1 0 5136 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3194
timestamp 1626908933
transform 1 0 5136 0 1 3885
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_610
timestamp 1626908933
transform 1 0 5280 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1332
timestamp 1626908933
transform 1 0 5280 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1092
timestamp 1626908933
transform 1 0 6048 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_494
timestamp 1626908933
transform 1 0 6048 0 1 3996
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1245
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_597
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1245
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_597
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1549
timestamp 1626908933
transform 1 0 6432 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_558
timestamp 1626908933
transform 1 0 6432 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1303
timestamp 1626908933
transform 1 0 6528 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_581
timestamp 1626908933
transform 1 0 6528 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_898
timestamp 1626908933
transform 1 0 7296 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_297
timestamp 1626908933
transform 1 0 7296 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1071
timestamp 1626908933
transform 1 0 7488 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_473
timestamp 1626908933
transform 1 0 7488 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1282
timestamp 1626908933
transform 1 0 7872 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_560
timestamp 1626908933
transform 1 0 7872 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3907
timestamp 1626908933
transform 1 0 8208 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1940
timestamp 1626908933
transform 1 0 8208 0 1 4403
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_450
timestamp 1626908933
transform 1 0 8640 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1048
timestamp 1626908933
transform 1 0 8640 0 1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_815
timestamp 1626908933
transform 1 0 8592 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2782
timestamp 1626908933
transform 1 0 8592 0 1 4329
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1221
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_573
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1221
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_573
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2787
timestamp 1626908933
transform 1 0 9168 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2784
timestamp 1626908933
transform 1 0 9072 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_852
timestamp 1626908933
transform 1 0 9168 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_849
timestamp 1626908933
transform 1 0 9072 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2784
timestamp 1626908933
transform 1 0 8784 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2778
timestamp 1626908933
transform 1 0 9168 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_817
timestamp 1626908933
transform 1 0 8784 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_811
timestamp 1626908933
transform 1 0 9168 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_88
timestamp 1626908933
transform 1 0 9024 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_26
timestamp 1626908933
transform 1 0 9024 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_439
timestamp 1626908933
transform 1 0 9408 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1037
timestamp 1626908933
transform 1 0 9408 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_557
timestamp 1626908933
transform 1 0 9312 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1548
timestamp 1626908933
transform 1 0 9312 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_846
timestamp 1626908933
transform 1 0 9264 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2781
timestamp 1626908933
transform 1 0 9264 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_556
timestamp 1626908933
transform 1 0 9792 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1547
timestamp 1626908933
transform 1 0 9792 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_128
timestamp 1626908933
transform 1 0 9744 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2095
timestamp 1626908933
transform 1 0 9744 0 1 3885
box -32 -32 32 32
use L1M1_PR  L1M1_PR_139
timestamp 1626908933
transform 1 0 9744 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2074
timestamp 1626908933
transform 1 0 9744 0 1 3885
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_305
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_662
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_694
timestamp 1626908933
transform 1 0 9888 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1685
timestamp 1626908933
transform 1 0 9888 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1560
timestamp 1626908933
transform 1 0 10128 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3495
timestamp 1626908933
transform 1 0 10128 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1726
timestamp 1626908933
transform 1 0 10320 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3693
timestamp 1626908933
transform 1 0 10320 0 1 4403
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1908
timestamp 1626908933
transform 1 0 10512 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3843
timestamp 1626908933
transform 1 0 10512 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_915
timestamp 1626908933
transform 1 0 10800 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2882
timestamp 1626908933
transform 1 0 10800 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1472
timestamp 1626908933
transform 1 0 10992 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3439
timestamp 1626908933
transform 1 0 10992 0 1 4255
box -32 -32 32 32
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_28
timestamp 1626908933
transform 1 0 10080 0 1 3996
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_4
timestamp 1626908933
transform 1 0 10080 0 1 3996
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1197
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_549
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1197
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_549
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1973
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_38
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2004
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_37
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1195
timestamp 1626908933
transform 1 0 12384 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_473
timestamp 1626908933
transform 1 0 12384 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_695
timestamp 1626908933
transform 1 0 13152 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1686
timestamp 1626908933
transform 1 0 13152 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_132
timestamp 1626908933
transform 1 0 12912 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_913
timestamp 1626908933
transform 1 0 13104 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2099
timestamp 1626908933
transform 1 0 12912 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2880
timestamp 1626908933
transform 1 0 13104 0 1 4477
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_32
timestamp 1626908933
transform 1 0 13248 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_93
timestamp 1626908933
transform 1 0 13248 0 1 3996
box -38 -49 326 715
use L1M1_PR  L1M1_PR_144
timestamp 1626908933
transform 1 0 13488 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_966
timestamp 1626908933
transform 1 0 13200 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_972
timestamp 1626908933
transform 1 0 13488 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2079
timestamp 1626908933
transform 1 0 13488 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2901
timestamp 1626908933
transform 1 0 13200 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2907
timestamp 1626908933
transform 1 0 13488 0 1 4107
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_448
timestamp 1626908933
transform 1 0 13536 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1170
timestamp 1626908933
transform 1 0 13536 0 1 3996
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1173
timestamp 1626908933
transform 1 0 13700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_525
timestamp 1626908933
transform 1 0 13700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1173
timestamp 1626908933
transform 1 0 13700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_525
timestamp 1626908933
transform 1 0 13700 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_919
timestamp 1626908933
transform 1 0 13872 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1935
timestamp 1626908933
transform 1 0 14640 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2886
timestamp 1626908933
transform 1 0 13872 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3902
timestamp 1626908933
transform 1 0 14640 0 1 3811
box -32 -32 32 32
use L1M1_PR  L1M1_PR_970
timestamp 1626908933
transform 1 0 14256 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1606
timestamp 1626908933
transform 1 0 14544 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2905
timestamp 1626908933
transform 1 0 14256 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3541
timestamp 1626908933
transform 1 0 14544 0 1 4107
box -29 -23 29 23
use M1M2_PR  M1M2_PR_925
timestamp 1626908933
transform 1 0 14256 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2892
timestamp 1626908933
transform 1 0 14256 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_722
timestamp 1626908933
transform 1 0 14448 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_976
timestamp 1626908933
transform 1 0 14640 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2657
timestamp 1626908933
transform 1 0 14448 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2911
timestamp 1626908933
transform 1 0 14640 0 1 4255
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_28
timestamp 1626908933
transform 1 0 14304 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_90
timestamp 1626908933
transform 1 0 14304 0 1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3485
timestamp 1626908933
transform 1 0 14832 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1518
timestamp 1626908933
transform 1 0 14832 0 1 4107
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1687
timestamp 1626908933
transform 1 0 14880 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_696
timestamp 1626908933
transform 1 0 14880 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_661
timestamp 1626908933
transform 1 0 14976 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_304
timestamp 1626908933
transform 1 0 14976 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_984
timestamp 1626908933
transform 1 0 15072 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_983
timestamp 1626908933
transform 1 0 14688 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_383
timestamp 1626908933
transform 1 0 15072 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_382
timestamp 1626908933
transform 1 0 14688 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_697
timestamp 1626908933
transform 1 0 15264 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1688
timestamp 1626908933
transform 1 0 15264 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_702
timestamp 1626908933
transform 1 0 15120 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2669
timestamp 1626908933
transform 1 0 15120 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_720
timestamp 1626908933
transform 1 0 15408 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2655
timestamp 1626908933
transform 1 0 15408 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_100
timestamp 1626908933
transform -1 0 15840 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_31
timestamp 1626908933
transform -1 0 15840 0 1 3996
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1149
timestamp 1626908933
transform 1 0 16100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_501
timestamp 1626908933
transform 1 0 16100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1149
timestamp 1626908933
transform 1 0 16100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_501
timestamp 1626908933
transform 1 0 16100 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2087
timestamp 1626908933
transform 1 0 15792 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_152
timestamp 1626908933
transform 1 0 15792 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1117
timestamp 1626908933
transform 1 0 15840 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_395
timestamp 1626908933
transform 1 0 15840 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2683
timestamp 1626908933
transform 1 0 16464 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_716
timestamp 1626908933
transform 1 0 16464 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2675
timestamp 1626908933
transform 1 0 16656 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2543
timestamp 1626908933
transform 1 0 16752 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_740
timestamp 1626908933
transform 1 0 16656 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_608
timestamp 1626908933
transform 1 0 16752 0 1 4551
box -29 -23 29 23
use M1M2_PR  M1M2_PR_138
timestamp 1626908933
transform 1 0 16848 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2105
timestamp 1626908933
transform 1 0 16848 0 1 3885
box -32 -32 32 32
use L1M1_PR  L1M1_PR_151
timestamp 1626908933
transform 1 0 16848 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2086
timestamp 1626908933
transform 1 0 16848 0 1 3885
box -29 -23 29 23
use M1M2_PR  M1M2_PR_137
timestamp 1626908933
transform 1 0 16848 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2104
timestamp 1626908933
transform 1 0 16848 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_150
timestamp 1626908933
transform 1 0 16848 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2085
timestamp 1626908933
transform 1 0 16848 0 1 4255
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_555
timestamp 1626908933
transform 1 0 16896 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1546
timestamp 1626908933
transform 1 0 16896 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_67
timestamp 1626908933
transform 1 0 16608 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_6
timestamp 1626908933
transform 1 0 16608 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_369
timestamp 1626908933
transform 1 0 16992 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1091
timestamp 1626908933
transform 1 0 16992 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1933
timestamp 1626908933
transform 1 0 18096 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3900
timestamp 1626908933
transform 1 0 18096 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_689
timestamp 1626908933
transform 1 0 18096 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2656
timestamp 1626908933
transform 1 0 18096 0 1 4477
box -32 -32 32 32
use L1M1_PR  L1M1_PR_209
timestamp 1626908933
transform 1 0 18192 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_706
timestamp 1626908933
transform 1 0 18096 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2144
timestamp 1626908933
transform 1 0 18192 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2641
timestamp 1626908933
transform 1 0 18096 0 1 4477
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_84
timestamp 1626908933
transform -1 0 18240 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_15
timestamp 1626908933
transform -1 0 18240 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_339
timestamp 1626908933
transform 1 0 18240 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1061
timestamp 1626908933
transform 1 0 18240 0 1 3996
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2143
timestamp 1626908933
transform 1 0 18576 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_208
timestamp 1626908933
transform 1 0 18576 0 1 3885
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1125
timestamp 1626908933
transform 1 0 18500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_477
timestamp 1626908933
transform 1 0 18500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1125
timestamp 1626908933
transform 1 0 18500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_477
timestamp 1626908933
transform 1 0 18500 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2864
timestamp 1626908933
transform 1 0 18288 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_897
timestamp 1626908933
transform 1 0 18288 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2567
timestamp 1626908933
transform 1 0 18288 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_600
timestamp 1626908933
transform 1 0 18288 0 1 4551
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_23
timestamp 1626908933
transform 1 0 19008 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_84
timestamp 1626908933
transform 1 0 19008 0 1 3996
box -38 -49 326 715
use M1M2_PR  M1M2_PR_188
timestamp 1626908933
transform 1 0 18672 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_189
timestamp 1626908933
transform 1 0 18672 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_976
timestamp 1626908933
transform 1 0 18864 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2155
timestamp 1626908933
transform 1 0 18672 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2156
timestamp 1626908933
transform 1 0 18672 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2943
timestamp 1626908933
transform 1 0 18864 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1039
timestamp 1626908933
transform 1 0 19056 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2974
timestamp 1626908933
transform 1 0 19056 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2880
timestamp 1626908933
transform 1 0 19248 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2142
timestamp 1626908933
transform 1 0 19248 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_945
timestamp 1626908933
transform 1 0 19248 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_207
timestamp 1626908933
transform 1 0 19248 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2863
timestamp 1626908933
transform 1 0 19248 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_896
timestamp 1626908933
transform 1 0 19248 0 1 4107
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_897
timestamp 1626908933
transform 1 0 19296 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_296
timestamp 1626908933
transform 1 0 19296 0 1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1932
timestamp 1626908933
transform 1 0 19440 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3899
timestamp 1626908933
transform 1 0 19440 0 1 3811
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2140
timestamp 1626908933
transform 1 0 19824 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_205
timestamp 1626908933
transform 1 0 19824 0 1 3885
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2154
timestamp 1626908933
transform 1 0 19824 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2153
timestamp 1626908933
transform 1 0 19824 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_187
timestamp 1626908933
transform 1 0 19824 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_186
timestamp 1626908933
transform 1 0 19824 0 1 4255
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1689
timestamp 1626908933
transform 1 0 19872 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_698
timestamp 1626908933
transform 1 0 19872 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1545
timestamp 1626908933
transform 1 0 20064 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_554
timestamp 1626908933
transform 1 0 20064 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_660
timestamp 1626908933
transform 1 0 19968 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_303
timestamp 1626908933
transform 1 0 19968 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_219
timestamp 1626908933
transform 1 0 20160 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_231
timestamp 1626908933
transform 1 0 19488 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_817
timestamp 1626908933
transform 1 0 20160 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_829
timestamp 1626908933
transform 1 0 19488 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_8
timestamp 1626908933
transform -1 0 20832 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_69
timestamp 1626908933
transform -1 0 20832 0 1 3996
box -38 -49 326 715
use M1M2_PR  M1M2_PR_692
timestamp 1626908933
transform 1 0 20400 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2659
timestamp 1626908933
transform 1 0 20400 0 1 4551
box -32 -32 32 32
use L1M1_PR  L1M1_PR_204
timestamp 1626908933
transform 1 0 20592 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2139
timestamp 1626908933
transform 1 0 20592 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_707
timestamp 1626908933
transform 1 0 20688 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_761
timestamp 1626908933
transform 1 0 20880 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2642
timestamp 1626908933
transform 1 0 20688 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2696
timestamp 1626908933
transform 1 0 20880 0 1 4107
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_453
timestamp 1626908933
transform 1 0 20900 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1101
timestamp 1626908933
transform 1 0 20900 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_453
timestamp 1626908933
transform 1 0 20900 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1101
timestamp 1626908933
transform 1 0 20900 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_0
timestamp 1626908933
transform 1 0 20832 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_23
timestamp 1626908933
transform 1 0 20832 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_736
timestamp 1626908933
transform 1 0 21072 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_795
timestamp 1626908933
transform 1 0 21456 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2703
timestamp 1626908933
transform 1 0 21072 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2762
timestamp 1626908933
transform 1 0 21456 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_794
timestamp 1626908933
transform 1 0 21456 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2761
timestamp 1626908933
transform 1 0 21456 0 1 4551
box -32 -32 32 32
use L1M1_PR  L1M1_PR_203
timestamp 1626908933
transform 1 0 21648 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_829
timestamp 1626908933
transform 1 0 21744 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2138
timestamp 1626908933
transform 1 0 21648 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2764
timestamp 1626908933
transform 1 0 21744 0 1 4551
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_108
timestamp 1626908933
transform 1 0 21600 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_39
timestamp 1626908933
transform 1 0 21600 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_785
timestamp 1626908933
transform 1 0 22080 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_187
timestamp 1626908933
transform 1 0 22080 0 1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2763
timestamp 1626908933
transform 1 0 22896 0 1 3811
box -29 -23 29 23
use L1M1_PR  L1M1_PR_828
timestamp 1626908933
transform 1 0 22896 0 1 3811
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1544
timestamp 1626908933
transform 1 0 22464 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_553
timestamp 1626908933
transform 1 0 22464 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_980
timestamp 1626908933
transform 1 0 22560 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_258
timestamp 1626908933
transform 1 0 22560 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_552
timestamp 1626908933
transform 1 0 23328 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1543
timestamp 1626908933
transform 1 0 23328 0 1 3996
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_429
timestamp 1626908933
transform 1 0 23300 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1077
timestamp 1626908933
transform 1 0 23300 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_429
timestamp 1626908933
transform 1 0 23300 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1077
timestamp 1626908933
transform 1 0 23300 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_100
timestamp 1626908933
transform 1 0 23664 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_573
timestamp 1626908933
transform 1 0 23472 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2067
timestamp 1626908933
transform 1 0 23664 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2540
timestamp 1626908933
transform 1 0 23472 0 1 4551
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_226
timestamp 1626908933
transform 1 0 23424 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_948
timestamp 1626908933
transform 1 0 23424 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_10
timestamp 1626908933
transform -1 0 24480 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_71
timestamp 1626908933
transform -1 0 24480 0 1 3996
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2513
timestamp 1626908933
transform 1 0 24336 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2049
timestamp 1626908933
transform 1 0 24240 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_578
timestamp 1626908933
transform 1 0 24336 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_114
timestamp 1626908933
transform 1 0 24240 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2682
timestamp 1626908933
transform 1 0 24432 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_747
timestamp 1626908933
transform 1 0 24432 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2690
timestamp 1626908933
transform 1 0 24528 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2689
timestamp 1626908933
transform 1 0 24528 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_723
timestamp 1626908933
transform 1 0 24528 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_722
timestamp 1626908933
transform 1 0 24528 0 1 4255
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1542
timestamp 1626908933
transform 1 0 24480 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_551
timestamp 1626908933
transform 1 0 24480 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_139
timestamp 1626908933
transform 1 0 24576 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_737
timestamp 1626908933
transform 1 0 24576 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_302
timestamp 1626908933
transform 1 0 24960 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_659
timestamp 1626908933
transform 1 0 24960 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_550
timestamp 1626908933
transform 1 0 25056 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1541
timestamp 1626908933
transform 1 0 25056 0 1 3996
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_405
timestamp 1626908933
transform 1 0 25700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1053
timestamp 1626908933
transform 1 0 25700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_405
timestamp 1626908933
transform 1 0 25700 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1053
timestamp 1626908933
transform 1 0 25700 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_194
timestamp 1626908933
transform 1 0 25152 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_916
timestamp 1626908933
transform 1 0 25152 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_295
timestamp 1626908933
transform 1 0 25920 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_896
timestamp 1626908933
transform 1 0 25920 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_549
timestamp 1626908933
transform 1 0 26112 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1540
timestamp 1626908933
transform 1 0 26112 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_970
timestamp 1626908933
transform 1 0 25968 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2937
timestamp 1626908933
transform 1 0 25968 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_745
timestamp 1626908933
transform 1 0 25776 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2680
timestamp 1626908933
transform 1 0 25776 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2969
timestamp 1626908933
transform 1 0 26256 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2137
timestamp 1626908933
transform 1 0 26160 0 1 3811
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1034
timestamp 1626908933
transform 1 0 26256 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_202
timestamp 1626908933
transform 1 0 26160 0 1 3811
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2152
timestamp 1626908933
transform 1 0 26160 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_185
timestamp 1626908933
transform 1 0 26160 0 1 3811
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2967
timestamp 1626908933
transform 1 0 26544 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2136
timestamp 1626908933
transform 1 0 26256 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1032
timestamp 1626908933
transform 1 0 26544 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_201
timestamp 1626908933
transform 1 0 26256 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2151
timestamp 1626908933
transform 1 0 26160 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_184
timestamp 1626908933
transform 1 0 26160 0 1 4255
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_85
timestamp 1626908933
transform -1 0 26496 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_24
timestamp 1626908933
transform -1 0 26496 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_1
timestamp 1626908933
transform 1 0 26496 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_24
timestamp 1626908933
transform 1 0 26496 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2936
timestamp 1626908933
transform 1 0 26640 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_969
timestamp 1626908933
transform 1 0 26640 0 1 4403
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_895
timestamp 1626908933
transform 1 0 27264 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_294
timestamp 1626908933
transform 1 0 27264 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_856
timestamp 1626908933
transform 1 0 27456 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_134
timestamp 1626908933
transform 1 0 27456 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1488
timestamp 1626908933
transform 1 0 28272 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3455
timestamp 1626908933
transform 1 0 28272 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1575
timestamp 1626908933
transform 1 0 28272 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3510
timestamp 1626908933
transform 1 0 28272 0 1 4107
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_381
timestamp 1626908933
transform 1 0 28100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1029
timestamp 1626908933
transform 1 0 28100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_381
timestamp 1626908933
transform 1 0 28100 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1029
timestamp 1626908933
transform 1 0 28100 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1033
timestamp 1626908933
transform 1 0 28464 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2968
timestamp 1626908933
transform 1 0 28464 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_22
timestamp 1626908933
transform 1 0 28224 0 1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_61
timestamp 1626908933
transform 1 0 28224 0 1 3996
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2964
timestamp 1626908933
transform 1 0 28656 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2135
timestamp 1626908933
transform 1 0 28752 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1029
timestamp 1626908933
transform 1 0 28656 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_200
timestamp 1626908933
transform 1 0 28752 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_894
timestamp 1626908933
transform 1 0 28800 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_293
timestamp 1626908933
transform 1 0 28800 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_821
timestamp 1626908933
transform 1 0 28992 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_99
timestamp 1626908933
transform 1 0 28992 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2149
timestamp 1626908933
transform 1 0 29616 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_182
timestamp 1626908933
transform 1 0 29616 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_893
timestamp 1626908933
transform 1 0 29760 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_892
timestamp 1626908933
transform 1 0 30048 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_292
timestamp 1626908933
transform 1 0 29760 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_291
timestamp 1626908933
transform 1 0 30048 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_658
timestamp 1626908933
transform 1 0 29952 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_301
timestamp 1626908933
transform 1 0 29952 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1539
timestamp 1626908933
transform 1 0 30240 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_548
timestamp 1626908933
transform 1 0 30240 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_784
timestamp 1626908933
transform 1 0 30336 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_62
timestamp 1626908933
transform 1 0 30336 0 1 3996
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1005
timestamp 1626908933
transform 1 0 30500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_357
timestamp 1626908933
transform 1 0 30500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1005
timestamp 1626908933
transform 1 0 30500 0 1 3996
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_357
timestamp 1626908933
transform 1 0 30500 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1538
timestamp 1626908933
transform 1 0 31104 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_547
timestamp 1626908933
transform 1 0 31104 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_742
timestamp 1626908933
transform 1 0 31200 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_20
timestamp 1626908933
transform 1 0 31200 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1690
timestamp 1626908933
transform 1 0 31968 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_699
timestamp 1626908933
transform 1 0 31968 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1699
timestamp 1626908933
transform 1 0 192 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_708
timestamp 1626908933
transform 1 0 192 0 1 5328
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_980
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_332
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_980
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_332
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1700
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_709
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_650
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_293
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_995
timestamp 1626908933
transform 1 0 0 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_891
timestamp 1626908933
transform 1 0 0 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_394
timestamp 1626908933
transform 1 0 0 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_290
timestamp 1626908933
transform 1 0 0 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_134
timestamp 1626908933
transform -1 0 960 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_65
timestamp 1626908933
transform -1 0 960 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_718
timestamp 1626908933
transform 1 0 192 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1440
timestamp 1626908933
transform 1 0 192 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_580
timestamp 1626908933
transform 1 0 960 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_581
timestamp 1626908933
transform 1 0 1056 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1178
timestamp 1626908933
transform 1 0 960 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1179
timestamp 1626908933
transform 1 0 1056 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_546
timestamp 1626908933
transform 1 0 960 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1537
timestamp 1626908933
transform 1 0 960 0 -1 5328
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_644
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1292
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_644
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1292
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__nor2_4  sky130_fd_sc_hs__nor2_4_1
timestamp 1626908933
transform 1 0 1344 0 1 5328
box -38 -49 902 715
use sky130_fd_sc_hs__nor2_4  sky130_fd_sc_hs__nor2_4_3
timestamp 1626908933
transform 1 0 1344 0 1 5328
box -38 -49 902 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_685
timestamp 1626908933
transform 1 0 1440 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1407
timestamp 1626908933
transform 1 0 1440 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_283
timestamp 1626908933
transform 1 0 2208 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_384
timestamp 1626908933
transform 1 0 2304 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_884
timestamp 1626908933
transform 1 0 2208 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_985
timestamp 1626908933
transform 1 0 2304 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_545
timestamp 1626908933
transform 1 0 2208 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1536
timestamp 1626908933
transform 1 0 2208 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1233
timestamp 1626908933
transform 1 0 2160 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3200
timestamp 1626908933
transform 1 0 2160 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3919
timestamp 1626908933
transform 1 0 2352 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1952
timestamp 1626908933
transform 1 0 2352 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_657
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_300
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3127
timestamp 1626908933
transform 1 0 2640 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1160
timestamp 1626908933
transform 1 0 2640 0 1 5143
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_986
timestamp 1626908933
transform 1 0 2592 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_385
timestamp 1626908933
transform 1 0 2592 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1149
timestamp 1626908933
transform 1 0 2400 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_551
timestamp 1626908933
transform 1 0 2400 0 1 5328
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_308
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_956
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_308
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_956
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1920
timestamp 1626908933
transform 1 0 2928 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3855
timestamp 1626908933
transform 1 0 2928 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_700
timestamp 1626908933
transform 1 0 2784 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_710
timestamp 1626908933
transform 1 0 2784 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1691
timestamp 1626908933
transform 1 0 2784 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1701
timestamp 1626908933
transform 1 0 2784 0 1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3249
timestamp 1626908933
transform 1 0 3216 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3165
timestamp 1626908933
transform 1 0 3024 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1314
timestamp 1626908933
transform 1 0 3216 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1230
timestamp 1626908933
transform 1 0 3024 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_883
timestamp 1626908933
transform 1 0 3168 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_282
timestamp 1626908933
transform 1 0 3168 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_117
timestamp 1626908933
transform 1 0 2880 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_56
timestamp 1626908933
transform 1 0 2880 0 1 5328
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3252
timestamp 1626908933
transform 1 0 3312 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3248
timestamp 1626908933
transform 1 0 3408 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1317
timestamp 1626908933
transform 1 0 3312 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1313
timestamp 1626908933
transform 1 0 3408 0 1 5143
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3201
timestamp 1626908933
transform 1 0 3312 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1234
timestamp 1626908933
transform 1 0 3312 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1137
timestamp 1626908933
transform 1 0 3456 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1136
timestamp 1626908933
transform 1 0 3360 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_539
timestamp 1626908933
transform 1 0 3456 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_538
timestamp 1626908933
transform 1 0 3360 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_10
timestamp 1626908933
transform -1 0 4224 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_2
timestamp 1626908933
transform -1 0 4224 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_5
timestamp 1626908933
transform 1 0 2880 0 -1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_11
timestamp 1626908933
transform 1 0 2880 0 -1 5328
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1268
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_620
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1268
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_620
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3198
timestamp 1626908933
transform 1 0 3888 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1231
timestamp 1626908933
transform 1 0 3888 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1692
timestamp 1626908933
transform 1 0 4032 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_701
timestamp 1626908933
transform 1 0 4032 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3245
timestamp 1626908933
transform 1 0 4176 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1310
timestamp 1626908933
transform 1 0 4176 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_996
timestamp 1626908933
transform 1 0 4224 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_987
timestamp 1626908933
transform 1 0 3840 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_395
timestamp 1626908933
transform 1 0 4224 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_386
timestamp 1626908933
transform 1 0 3840 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_521
timestamp 1626908933
transform 1 0 4608 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1119
timestamp 1626908933
transform 1 0 4608 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_711
timestamp 1626908933
transform 1 0 4416 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1702
timestamp 1626908933
transform 1 0 4416 0 1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1300
timestamp 1626908933
transform 1 0 4464 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1312
timestamp 1626908933
transform 1 0 4560 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3235
timestamp 1626908933
transform 1 0 4464 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3247
timestamp 1626908933
transform 1 0 4560 0 1 5069
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_130
timestamp 1626908933
transform 1 0 4512 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_61
timestamp 1626908933
transform 1 0 4512 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nor2_2  sky130_fd_sc_hs__nor2_2_0
timestamp 1626908933
transform -1 0 4608 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nor2_2  sky130_fd_sc_hs__nor2_2_2
timestamp 1626908933
transform -1 0 4608 0 -1 5328
box -38 -49 518 715
use M1M2_PR  M1M2_PR_3191
timestamp 1626908933
transform 1 0 4848 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1224
timestamp 1626908933
transform 1 0 4848 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_649
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_292
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_932
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_284
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_932
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_284
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3238
timestamp 1626908933
transform 1 0 5232 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1303
timestamp 1626908933
transform 1 0 5232 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3193
timestamp 1626908933
transform 1 0 5136 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1226
timestamp 1626908933
transform 1 0 5136 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_988
timestamp 1626908933
transform 1 0 4992 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_387
timestamp 1626908933
transform 1 0 4992 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1104
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_506
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1301
timestamp 1626908933
transform 1 0 5520 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3236
timestamp 1626908933
transform 1 0 5520 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_136
timestamp 1626908933
transform 1 0 5472 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_67
timestamp 1626908933
transform 1 0 5472 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nand4_2  sky130_fd_sc_hs__nand4_2_0
timestamp 1626908933
transform 1 0 5184 0 -1 5328
box -38 -49 998 715
use sky130_fd_sc_hs__nand4_2  sky130_fd_sc_hs__nand4_2_1
timestamp 1626908933
transform 1 0 5184 0 -1 5328
box -38 -49 998 715
use M1M2_PR  M1M2_PR_1155
timestamp 1626908933
transform 1 0 5808 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3122
timestamp 1626908933
transform 1 0 5808 0 1 5143
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1224
timestamp 1626908933
transform 1 0 6000 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1298
timestamp 1626908933
transform 1 0 5808 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1299
timestamp 1626908933
transform 1 0 6000 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3159
timestamp 1626908933
transform 1 0 6000 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3233
timestamp 1626908933
transform 1 0 5808 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3234
timestamp 1626908933
transform 1 0 6000 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_396
timestamp 1626908933
transform 1 0 5952 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_997
timestamp 1626908933
transform 1 0 5952 0 1 5328
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1222
timestamp 1626908933
transform 1 0 6672 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3189
timestamp 1626908933
transform 1 0 6672 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_13
timestamp 1626908933
transform 1 0 6912 0 -1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_52
timestamp 1626908933
transform 1 0 6912 0 -1 5328
box -38 -49 614 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_596
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1244
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_596
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1244
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_580
timestamp 1626908933
transform 1 0 6144 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1302
timestamp 1626908933
transform 1 0 6144 0 -1 5328
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3547
timestamp 1626908933
transform 1 0 6960 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1612
timestamp 1626908933
transform 1 0 6960 0 1 4773
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3491
timestamp 1626908933
transform 1 0 6960 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2877
timestamp 1626908933
transform 1 0 7056 0 1 4921
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1524
timestamp 1626908933
transform 1 0 6960 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_910
timestamp 1626908933
transform 1 0 7056 0 1 4921
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2900
timestamp 1626908933
transform 1 0 7152 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_965
timestamp 1626908933
transform 1 0 7152 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2896
timestamp 1626908933
transform 1 0 7344 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_961
timestamp 1626908933
transform 1 0 7344 0 1 4921
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_656
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_299
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_140
timestamp 1626908933
transform 1 0 7632 0 1 4847
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2075
timestamp 1626908933
transform 1 0 7632 0 1 4847
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_260
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_908
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_260
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_908
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_2
timestamp 1626908933
transform 1 0 7584 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_25
timestamp 1626908933
transform 1 0 7584 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_27
timestamp 1626908933
transform -1 0 8352 0 1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_2
timestamp 1626908933
transform -1 0 8352 0 1 5328
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_2783
timestamp 1626908933
transform 1 0 8304 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_848
timestamp 1626908933
transform 1 0 8304 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2786
timestamp 1626908933
transform 1 0 8496 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_851
timestamp 1626908933
transform 1 0 8496 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2781
timestamp 1626908933
transform 1 0 8592 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_814
timestamp 1626908933
transform 1 0 8592 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3498
timestamp 1626908933
transform 1 0 8592 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1563
timestamp 1626908933
transform 1 0 8592 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2790
timestamp 1626908933
transform 1 0 8688 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_855
timestamp 1626908933
transform 1 0 8688 0 1 5069
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3444
timestamp 1626908933
transform 1 0 8688 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1477
timestamp 1626908933
transform 1 0 8688 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_816
timestamp 1626908933
transform 1 0 8784 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2783
timestamp 1626908933
transform 1 0 8784 0 1 5069
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_572
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1220
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_572
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1220
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_544
timestamp 1626908933
transform 1 0 8736 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_712
timestamp 1626908933
transform 1 0 8736 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1535
timestamp 1626908933
transform 1 0 8736 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1703
timestamp 1626908933
transform 1 0 8736 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_86
timestamp 1626908933
transform -1 0 9312 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_17
timestamp 1626908933
transform -1 0 9312 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_540
timestamp 1626908933
transform 1 0 8832 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1262
timestamp 1626908933
transform 1 0 8832 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_455
timestamp 1626908933
transform 1 0 8352 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1053
timestamp 1626908933
transform 1 0 8352 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_14
timestamp 1626908933
transform 1 0 8352 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_76
timestamp 1626908933
transform 1 0 8352 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_537
timestamp 1626908933
transform 1 0 9312 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1528
timestamp 1626908933
transform 1 0 9312 0 1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_810
timestamp 1626908933
transform 1 0 9168 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2777
timestamp 1626908933
transform 1 0 9168 0 1 4773
box -32 -32 32 32
use L1M1_PR  L1M1_PR_958
timestamp 1626908933
transform 1 0 9552 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2893
timestamp 1626908933
transform 1 0 9552 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2899
timestamp 1626908933
transform 1 0 9744 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_964
timestamp 1626908933
transform 1 0 9744 0 1 5143
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2094
timestamp 1626908933
transform 1 0 9744 0 1 4847
box -32 -32 32 32
use M1M2_PR  M1M2_PR_127
timestamp 1626908933
transform 1 0 9744 0 1 4847
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2073
timestamp 1626908933
transform 1 0 9936 0 1 4847
box -29 -23 29 23
use L1M1_PR  L1M1_PR_138
timestamp 1626908933
transform 1 0 9936 0 1 4847
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1704
timestamp 1626908933
transform 1 0 9888 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1527
timestamp 1626908933
transform 1 0 9792 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_713
timestamp 1626908933
transform 1 0 9888 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_536
timestamp 1626908933
transform 1 0 9792 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_648
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_291
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_890
timestamp 1626908933
transform 1 0 9888 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_289
timestamp 1626908933
transform 1 0 9888 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_94
timestamp 1626908933
transform 1 0 9600 0 -1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_33
timestamp 1626908933
transform 1 0 9600 0 -1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_438
timestamp 1626908933
transform 1 0 9408 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1036
timestamp 1626908933
transform 1 0 9408 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_397
timestamp 1626908933
transform 1 0 10080 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_998
timestamp 1626908933
transform 1 0 10080 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_37
timestamp 1626908933
transform -1 0 10560 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_99
timestamp 1626908933
transform -1 0 10560 0 1 5328
box -38 -49 326 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_236
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_884
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_236
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_884
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2879
timestamp 1626908933
transform 1 0 10416 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_912
timestamp 1626908933
transform 1 0 10416 0 1 5143
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1526
timestamp 1626908933
transform 1 0 10560 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_535
timestamp 1626908933
transform 1 0 10560 0 1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2884
timestamp 1626908933
transform 1 0 10704 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2586
timestamp 1626908933
transform 1 0 10608 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_917
timestamp 1626908933
transform 1 0 10704 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_619
timestamp 1626908933
transform 1 0 10608 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2897
timestamp 1626908933
transform 1 0 10800 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_962
timestamp 1626908933
transform 1 0 10800 0 1 5143
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_497
timestamp 1626908933
transform 1 0 10656 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_521
timestamp 1626908933
transform 1 0 10080 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1219
timestamp 1626908933
transform 1 0 10656 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1243
timestamp 1626908933
transform 1 0 10080 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_89
timestamp 1626908933
transform 1 0 10848 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_27
timestamp 1626908933
transform 1 0 10848 0 -1 5328
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2562
timestamp 1626908933
transform 1 0 10992 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_627
timestamp 1626908933
transform 1 0 10992 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2730
timestamp 1626908933
transform 1 0 10896 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_763
timestamp 1626908933
transform 1 0 10896 0 1 4773
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2903
timestamp 1626908933
transform 1 0 11184 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_968
timestamp 1626908933
transform 1 0 11184 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3544
timestamp 1626908933
transform 1 0 11088 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1609
timestamp 1626908933
transform 1 0 11088 0 1 5217
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3490
timestamp 1626908933
transform 1 0 11088 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1523
timestamp 1626908933
transform 1 0 11088 0 1 5217
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1196
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_548
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1196
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_548
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_543
timestamp 1626908933
transform 1 0 11232 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1534
timestamp 1626908933
transform 1 0 11232 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_792
timestamp 1626908933
transform 1 0 11856 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2727
timestamp 1626908933
transform 1 0 11856 0 1 4773
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_87
timestamp 1626908933
transform -1 0 12192 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_18
timestamp 1626908933
transform -1 0 12192 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_400
timestamp 1626908933
transform 1 0 11328 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_998
timestamp 1626908933
transform 1 0 11328 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_1
timestamp 1626908933
transform -1 0 12000 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_7
timestamp 1626908933
transform -1 0 12000 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_281
timestamp 1626908933
transform 1 0 12000 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_388
timestamp 1626908933
transform 1 0 12192 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_882
timestamp 1626908933
transform 1 0 12000 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_989
timestamp 1626908933
transform 1 0 12192 0 -1 5328
box -38 -49 230 715
use L1M1_PR  L1M1_PR_39
timestamp 1626908933
transform 1 0 12144 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1974
timestamp 1626908933
transform 1 0 12144 0 1 4995
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_212
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_860
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_212
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_860
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use M1M2_PR  M1M2_PR_36
timestamp 1626908933
transform 1 0 12336 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2003
timestamp 1626908933
transform 1 0 12336 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_298
timestamp 1626908933
transform 1 0 12480 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_655
timestamp 1626908933
transform 1 0 12480 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_702
timestamp 1626908933
transform 1 0 12384 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1693
timestamp 1626908933
transform 1 0 12384 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_74
timestamp 1626908933
transform 1 0 12576 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_5
timestamp 1626908933
transform 1 0 12576 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_472
timestamp 1626908933
transform 1 0 12192 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1194
timestamp 1626908933
transform 1 0 12192 0 1 5328
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2565
timestamp 1626908933
transform 1 0 12912 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1978
timestamp 1626908933
transform 1 0 12912 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_630
timestamp 1626908933
transform 1 0 12912 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_43
timestamp 1626908933
transform 1 0 12912 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2588
timestamp 1626908933
transform 1 0 12912 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2100
timestamp 1626908933
transform 1 0 12816 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_621
timestamp 1626908933
transform 1 0 12912 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_133
timestamp 1626908933
transform 1 0 12816 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_63
timestamp 1626908933
transform -1 0 13248 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_1
timestamp 1626908933
transform -1 0 13248 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_990
timestamp 1626908933
transform 1 0 13056 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_389
timestamp 1626908933
transform 1 0 13056 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_703
timestamp 1626908933
transform 1 0 13248 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1694
timestamp 1626908933
transform 1 0 13248 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_38
timestamp 1626908933
transform 1 0 13488 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2005
timestamp 1626908933
transform 1 0 13488 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_41
timestamp 1626908933
transform 1 0 13584 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_145
timestamp 1626908933
transform 1 0 13392 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1976
timestamp 1626908933
transform 1 0 13584 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2080
timestamp 1626908933
transform 1 0 13392 0 1 5069
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_4
timestamp 1626908933
transform 1 0 13248 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_27
timestamp 1626908933
transform 1 0 13248 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_3
timestamp 1626908933
transform 1 0 13344 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_28
timestamp 1626908933
transform 1 0 13344 0 -1 5328
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1172
timestamp 1626908933
transform 1 0 13700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_524
timestamp 1626908933
transform 1 0 13700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1172
timestamp 1626908933
transform 1 0 13700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_524
timestamp 1626908933
transform 1 0 13700 0 1 5328
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2551
timestamp 1626908933
transform 1 0 13680 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_616
timestamp 1626908933
transform 1 0 13680 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1533
timestamp 1626908933
transform 1 0 13824 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_542
timestamp 1626908933
transform 1 0 13824 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_346
timestamp 1626908933
transform 1 0 13920 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_944
timestamp 1626908933
transform 1 0 13920 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_13
timestamp 1626908933
transform 1 0 14304 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_65
timestamp 1626908933
transform 1 0 14304 0 1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_607
timestamp 1626908933
transform 1 0 14064 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2574
timestamp 1626908933
transform 1 0 14064 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_36
timestamp 1626908933
transform -1 0 14304 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_98
timestamp 1626908933
transform -1 0 14304 0 1 5328
box -38 -49 326 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_836
timestamp 1626908933
transform 1 0 14900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_188
timestamp 1626908933
transform 1 0 14900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_836
timestamp 1626908933
transform 1 0 14900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_188
timestamp 1626908933
transform 1 0 14900 0 1 4662
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3904
timestamp 1626908933
transform 1 0 14544 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1937
timestamp 1626908933
transform 1 0 14544 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_999
timestamp 1626908933
transform 1 0 14688 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_398
timestamp 1626908933
transform 1 0 14688 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1706
timestamp 1626908933
transform 1 0 15072 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1705
timestamp 1626908933
transform 1 0 14880 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1532
timestamp 1626908933
transform 1 0 15072 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_715
timestamp 1626908933
transform 1 0 15072 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_714
timestamp 1626908933
transform 1 0 14880 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_541
timestamp 1626908933
transform 1 0 15072 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_647
timestamp 1626908933
transform 1 0 14976 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_290
timestamp 1626908933
transform 1 0 14976 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_65
timestamp 1626908933
transform 1 0 15168 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_4
timestamp 1626908933
transform 1 0 15168 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_433
timestamp 1626908933
transform 1 0 14304 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1155
timestamp 1626908933
transform 1 0 14304 0 -1 5328
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1554
timestamp 1626908933
transform 1 0 15216 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1902
timestamp 1626908933
transform 1 0 15600 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3489
timestamp 1626908933
transform 1 0 15216 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3837
timestamp 1626908933
transform 1 0 15600 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1469
timestamp 1626908933
transform 1 0 16272 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3436
timestamp 1626908933
transform 1 0 16272 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_3
timestamp 1626908933
transform 1 0 16224 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_42
timestamp 1626908933
transform 1 0 16224 0 1 5328
box -38 -49 614 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_500
timestamp 1626908933
transform 1 0 16100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1148
timestamp 1626908933
transform 1 0 16100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_500
timestamp 1626908933
transform 1 0 16100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1148
timestamp 1626908933
transform 1 0 16100 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_415
timestamp 1626908933
transform 1 0 15456 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1137
timestamp 1626908933
transform 1 0 15456 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_31
timestamp 1626908933
transform 1 0 15168 0 -1 5328
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_7
timestamp 1626908933
transform 1 0 15168 0 -1 5328
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_45
timestamp 1626908933
transform 1 0 16752 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2012
timestamp 1626908933
transform 1 0 16752 0 1 5217
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_164
timestamp 1626908933
transform 1 0 17300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_812
timestamp 1626908933
transform 1 0 17300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_164
timestamp 1626908933
transform 1 0 17300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_812
timestamp 1626908933
transform 1 0 17300 0 1 4662
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1704
timestamp 1626908933
transform 1 0 17328 0 1 4921
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3671
timestamp 1626908933
transform 1 0 17328 0 1 4921
box -32 -32 32 32
use L1M1_PR  L1M1_PR_49
timestamp 1626908933
transform 1 0 17424 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1984
timestamp 1626908933
transform 1 0 17424 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_297
timestamp 1626908933
transform 1 0 17472 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_654
timestamp 1626908933
transform 1 0 17472 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_540
timestamp 1626908933
transform 1 0 17568 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_716
timestamp 1626908933
transform 1 0 17568 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1531
timestamp 1626908933
transform 1 0 17568 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1707
timestamp 1626908933
transform 1 0 17568 0 1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2162
timestamp 1626908933
transform 1 0 17712 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_195
timestamp 1626908933
transform 1 0 17712 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_871
timestamp 1626908933
transform 1 0 17664 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_273
timestamp 1626908933
transform 1 0 17664 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_386
timestamp 1626908933
transform 1 0 16800 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1108
timestamp 1626908933
transform 1 0 16800 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_539
timestamp 1626908933
transform 1 0 18048 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1530
timestamp 1626908933
transform 1 0 18048 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_688
timestamp 1626908933
transform 1 0 18096 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2655
timestamp 1626908933
transform 1 0 18096 0 1 4773
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_476
timestamp 1626908933
transform 1 0 18500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1124
timestamp 1626908933
transform 1 0 18500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_476
timestamp 1626908933
transform 1 0 18500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1124
timestamp 1626908933
transform 1 0 18500 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1695
timestamp 1626908933
transform 1 0 18912 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_704
timestamp 1626908933
transform 1 0 18912 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2879
timestamp 1626908933
transform 1 0 19344 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2146
timestamp 1626908933
transform 1 0 19344 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_944
timestamp 1626908933
transform 1 0 19344 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_211
timestamp 1626908933
transform 1 0 19344 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2862
timestamp 1626908933
transform 1 0 19248 0 1 4921
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2160
timestamp 1626908933
transform 1 0 19248 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_895
timestamp 1626908933
transform 1 0 19248 0 1 4921
box -32 -32 32 32
use M1M2_PR  M1M2_PR_193
timestamp 1626908933
transform 1 0 19248 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_362
timestamp 1626908933
transform 1 0 18144 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1084
timestamp 1626908933
transform 1 0 18144 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_1
timestamp 1626908933
transform 1 0 19008 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_9
timestamp 1626908933
transform 1 0 19008 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_49
timestamp 1626908933
transform -1 0 19872 0 1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_24
timestamp 1626908933
transform -1 0 19872 0 1 5328
box -38 -49 2246 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_788
timestamp 1626908933
transform 1 0 19700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_140
timestamp 1626908933
transform 1 0 19700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_788
timestamp 1626908933
transform 1 0 19700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_140
timestamp 1626908933
transform 1 0 19700 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3505
timestamp 1626908933
transform 1 0 19632 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1570
timestamp 1626908933
transform 1 0 19632 0 1 5217
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3450
timestamp 1626908933
transform 1 0 19728 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1483
timestamp 1626908933
transform 1 0 19728 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1708
timestamp 1626908933
transform 1 0 19872 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_717
timestamp 1626908933
transform 1 0 19872 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_646
timestamp 1626908933
transform 1 0 19968 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_289
timestamp 1626908933
transform 1 0 19968 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_822
timestamp 1626908933
transform 1 0 19680 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_224
timestamp 1626908933
transform 1 0 19680 0 -1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_111
timestamp 1626908933
transform 1 0 20112 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2078
timestamp 1626908933
transform 1 0 20112 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_310
timestamp 1626908933
transform 1 0 20064 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1032
timestamp 1626908933
transform 1 0 20064 0 -1 5328
box -38 -49 806 715
use L1M1_PR  L1M1_PR_703
timestamp 1626908933
transform 1 0 20784 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2638
timestamp 1626908933
transform 1 0 20784 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_120
timestamp 1626908933
transform 1 0 21072 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2055
timestamp 1626908933
transform 1 0 21072 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_570
timestamp 1626908933
transform 1 0 21072 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2537
timestamp 1626908933
transform 1 0 21072 0 1 5217
box -32 -32 32 32
use L1M1_PR  L1M1_PR_574
timestamp 1626908933
transform 1 0 21072 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2509
timestamp 1626908933
transform 1 0 21072 0 1 5217
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_452
timestamp 1626908933
transform 1 0 20900 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1100
timestamp 1626908933
transform 1 0 20900 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_452
timestamp 1626908933
transform 1 0 20900 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1100
timestamp 1626908933
transform 1 0 20900 0 1 5328
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2765
timestamp 1626908933
transform 1 0 21360 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2053
timestamp 1626908933
transform 1 0 21168 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_830
timestamp 1626908933
transform 1 0 21360 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_118
timestamp 1626908933
transform 1 0 21168 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2071
timestamp 1626908933
transform 1 0 21168 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_104
timestamp 1626908933
transform 1 0 21168 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_889
timestamp 1626908933
transform 1 0 21408 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_288
timestamp 1626908933
transform 1 0 21408 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_16
timestamp 1626908933
transform 1 0 20832 0 -1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_3
timestamp 1626908933
transform 1 0 20832 0 -1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_538
timestamp 1626908933
transform 1 0 21600 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1529
timestamp 1626908933
transform 1 0 21600 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_793
timestamp 1626908933
transform 1 0 21456 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2760
timestamp 1626908933
transform 1 0 21456 0 1 4995
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_116
timestamp 1626908933
transform 1 0 22100 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_764
timestamp 1626908933
transform 1 0 22100 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_116
timestamp 1626908933
transform 1 0 22100 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_764
timestamp 1626908933
transform 1 0 22100 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_274
timestamp 1626908933
transform 1 0 21696 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_996
timestamp 1626908933
transform 1 0 21696 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_46
timestamp 1626908933
transform -1 0 22368 0 1 5328
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_22
timestamp 1626908933
transform -1 0 22368 0 1 5328
box -38 -49 2342 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1000
timestamp 1626908933
transform 1 0 22368 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_399
timestamp 1626908933
transform 1 0 22368 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1709
timestamp 1626908933
transform 1 0 22560 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_718
timestamp 1626908933
transform 1 0 22560 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_991
timestamp 1626908933
transform 1 0 22560 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_390
timestamp 1626908933
transform 1 0 22560 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_653
timestamp 1626908933
transform 1 0 22464 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_296
timestamp 1626908933
transform 1 0 22464 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3410
timestamp 1626908933
transform 1 0 22800 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1443
timestamp 1626908933
transform 1 0 22800 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1696
timestamp 1626908933
transform 1 0 22752 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_705
timestamp 1626908933
transform 1 0 22752 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_935
timestamp 1626908933
transform 1 0 22896 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2870
timestamp 1626908933
transform 1 0 22896 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_826
timestamp 1626908933
transform 1 0 23088 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2761
timestamp 1626908933
transform 1 0 23088 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1527
timestamp 1626908933
transform 1 0 22992 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3462
timestamp 1626908933
transform 1 0 22992 0 1 5217
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_428
timestamp 1626908933
transform 1 0 23300 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1076
timestamp 1626908933
transform 1 0 23300 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_428
timestamp 1626908933
transform 1 0 23300 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1076
timestamp 1626908933
transform 1 0 23300 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_85
timestamp 1626908933
transform -1 0 23232 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_23
timestamp 1626908933
transform -1 0 23232 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_3
timestamp 1626908933
transform 1 0 23232 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_26
timestamp 1626908933
transform 1 0 23232 0 -1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_792
timestamp 1626908933
transform 1 0 23760 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_884
timestamp 1626908933
transform 1 0 23664 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2759
timestamp 1626908933
transform 1 0 23760 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2851
timestamp 1626908933
transform 1 0 23664 0 1 5143
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1697
timestamp 1626908933
transform 1 0 24192 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_706
timestamp 1626908933
transform 1 0 24192 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2866
timestamp 1626908933
transform 1 0 24240 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_931
timestamp 1626908933
transform 1 0 24240 0 1 5217
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2850
timestamp 1626908933
transform 1 0 24240 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_883
timestamp 1626908933
transform 1 0 24240 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_79
timestamp 1626908933
transform -1 0 24576 0 -1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_17
timestamp 1626908933
transform -1 0 24576 0 -1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_992
timestamp 1626908933
transform 1 0 24000 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_391
timestamp 1626908933
transform 1 0 24000 0 -1 5328
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_740
timestamp 1626908933
transform 1 0 24500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_92
timestamp 1626908933
transform 1 0 24500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_740
timestamp 1626908933
transform 1 0 24500 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_92
timestamp 1626908933
transform 1 0 24500 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2867
timestamp 1626908933
transform 1 0 24432 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2759
timestamp 1626908933
transform 1 0 24528 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_932
timestamp 1626908933
transform 1 0 24432 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_824
timestamp 1626908933
transform 1 0 24528 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_888
timestamp 1626908933
transform 1 0 24576 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_287
timestamp 1626908933
transform 1 0 24576 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_736
timestamp 1626908933
transform 1 0 24768 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_138
timestamp 1626908933
transform 1 0 24768 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_43
timestamp 1626908933
transform 1 0 22656 0 1 5328
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_19
timestamp 1626908933
transform 1 0 22656 0 1 5328
box -38 -49 2342 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_288
timestamp 1626908933
transform 1 0 24960 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_645
timestamp 1626908933
transform 1 0 24960 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_534
timestamp 1626908933
transform 1 0 25056 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1525
timestamp 1626908933
transform 1 0 25056 0 1 5328
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1052
timestamp 1626908933
transform 1 0 25700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_404
timestamp 1626908933
transform 1 0 25700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1052
timestamp 1626908933
transform 1 0 25700 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_404
timestamp 1626908933
transform 1 0 25700 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1524
timestamp 1626908933
transform 1 0 25920 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_533
timestamp 1626908933
transform 1 0 25920 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_887
timestamp 1626908933
transform 1 0 25920 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_286
timestamp 1626908933
transform 1 0 25920 0 -1 5328
box -38 -49 230 715
use M1M2_PR  M1M2_PR_2148
timestamp 1626908933
transform 1 0 26256 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_181
timestamp 1626908933
transform 1 0 26256 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_709
timestamp 1626908933
transform 1 0 26112 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_708
timestamp 1626908933
transform 1 0 26016 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_111
timestamp 1626908933
transform 1 0 26112 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_110
timestamp 1626908933
transform 1 0 26016 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_192
timestamp 1626908933
transform 1 0 25152 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_193
timestamp 1626908933
transform 1 0 25152 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_914
timestamp 1626908933
transform 1 0 25152 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_915
timestamp 1626908933
transform 1 0 25152 0 -1 5328
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_716
timestamp 1626908933
transform 1 0 26900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_68
timestamp 1626908933
transform 1 0 26900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_716
timestamp 1626908933
transform 1 0 26900 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_68
timestamp 1626908933
transform 1 0 26900 0 1 4662
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3458
timestamp 1626908933
transform 1 0 26736 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1491
timestamp 1626908933
transform 1 0 26736 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_881
timestamp 1626908933
transform 1 0 26784 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_280
timestamp 1626908933
transform 1 0 26784 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_97
timestamp 1626908933
transform 1 0 26400 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_35
timestamp 1626908933
transform 1 0 26400 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_295
timestamp 1626908933
transform 1 0 27456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_652
timestamp 1626908933
transform 1 0 27456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_392
timestamp 1626908933
transform 1 0 27264 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_993
timestamp 1626908933
transform 1 0 27264 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_532
timestamp 1626908933
transform 1 0 26976 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1523
timestamp 1626908933
transform 1 0 26976 0 1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1577
timestamp 1626908933
transform 1 0 27600 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3512
timestamp 1626908933
transform 1 0 27600 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_143
timestamp 1626908933
transform 1 0 27072 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_165
timestamp 1626908933
transform 1 0 26496 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_865
timestamp 1626908933
transform 1 0 27072 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_887
timestamp 1626908933
transform 1 0 26496 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_45
timestamp 1626908933
transform 1 0 27552 0 -1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_20
timestamp 1626908933
transform 1 0 27552 0 -1 5328
box -38 -49 2246 715
use M1M2_PR  M1M2_PR_1682
timestamp 1626908933
transform 1 0 27696 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3649
timestamp 1626908933
transform 1 0 27696 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1921
timestamp 1626908933
transform 1 0 27888 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3888
timestamp 1626908933
transform 1 0 27888 0 1 5069
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1890
timestamp 1626908933
transform 1 0 27888 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3825
timestamp 1626908933
transform 1 0 27888 0 1 5069
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_380
timestamp 1626908933
transform 1 0 28100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1028
timestamp 1626908933
transform 1 0 28100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_380
timestamp 1626908933
transform 1 0 28100 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1028
timestamp 1626908933
transform 1 0 28100 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_880
timestamp 1626908933
transform 1 0 27840 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_279
timestamp 1626908933
transform 1 0 27840 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_110
timestamp 1626908933
transform 1 0 28416 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_832
timestamp 1626908933
transform 1 0 28416 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_75
timestamp 1626908933
transform 1 0 28032 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_673
timestamp 1626908933
transform 1 0 28032 0 1 5328
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_692
timestamp 1626908933
transform 1 0 29300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_44
timestamp 1626908933
transform 1 0 29300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_692
timestamp 1626908933
transform 1 0 29300 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_44
timestamp 1626908933
transform 1 0 29300 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_798
timestamp 1626908933
transform 1 0 29184 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_76
timestamp 1626908933
transform 1 0 29184 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_285
timestamp 1626908933
transform 1 0 29760 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_886
timestamp 1626908933
transform 1 0 29760 0 -1 5328
box -38 -49 230 715
use L1M1_PR  L1M1_PR_196
timestamp 1626908933
transform 1 0 29712 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2131
timestamp 1626908933
transform 1 0 29712 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_287
timestamp 1626908933
transform 1 0 29952 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_644
timestamp 1626908933
transform 1 0 29952 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_278
timestamp 1626908933
transform 1 0 30048 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_879
timestamp 1626908933
transform 1 0 30048 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_35
timestamp 1626908933
transform 1 0 29952 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_633
timestamp 1626908933
transform 1 0 29952 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1522
timestamp 1626908933
transform 1 0 30240 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_531
timestamp 1626908933
transform 1 0 30240 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_783
timestamp 1626908933
transform 1 0 30336 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_782
timestamp 1626908933
transform 1 0 30336 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_61
timestamp 1626908933
transform 1 0 30336 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_60
timestamp 1626908933
transform 1 0 30336 0 1 5328
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_356
timestamp 1626908933
transform 1 0 30500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1004
timestamp 1626908933
transform 1 0 30500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_356
timestamp 1626908933
transform 1 0 30500 0 1 5328
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1004
timestamp 1626908933
transform 1 0 30500 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_530
timestamp 1626908933
transform 1 0 31104 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1521
timestamp 1626908933
transform 1 0 31104 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_19
timestamp 1626908933
transform 1 0 31200 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_741
timestamp 1626908933
transform 1 0 31200 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_13
timestamp 1626908933
transform 1 0 31104 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_611
timestamp 1626908933
transform 1 0 31104 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_284
timestamp 1626908933
transform 1 0 31488 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_885
timestamp 1626908933
transform 1 0 31488 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_294
timestamp 1626908933
transform 1 0 31680 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_651
timestamp 1626908933
transform 1 0 31680 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_393
timestamp 1626908933
transform 1 0 31776 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_994
timestamp 1626908933
transform 1 0 31776 0 -1 5328
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_20
timestamp 1626908933
transform 1 0 31700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_668
timestamp 1626908933
transform 1 0 31700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_20
timestamp 1626908933
transform 1 0 31700 0 1 4662
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_668
timestamp 1626908933
transform 1 0 31700 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_707
timestamp 1626908933
transform 1 0 31968 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_719
timestamp 1626908933
transform 1 0 31968 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1698
timestamp 1626908933
transform 1 0 31968 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1710
timestamp 1626908933
transform 1 0 31968 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_277
timestamp 1626908933
transform 1 0 0 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_878
timestamp 1626908933
transform 1 0 0 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1953
timestamp 1626908933
transform 1 0 144 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3920
timestamp 1626908933
transform 1 0 144 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3857
timestamp 1626908933
transform 1 0 624 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1922
timestamp 1626908933
transform 1 0 624 0 1 5661
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_979
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_331
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_979
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_331
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3281
timestamp 1626908933
transform 1 0 624 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1346
timestamp 1626908933
transform 1 0 624 0 1 5883
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3228
timestamp 1626908933
transform 1 0 720 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1261
timestamp 1626908933
transform 1 0 720 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_717
timestamp 1626908933
transform 1 0 192 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1439
timestamp 1626908933
transform 1 0 192 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_529
timestamp 1626908933
transform 1 0 960 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1520
timestamp 1626908933
transform 1 0 960 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1246
timestamp 1626908933
transform 1 0 1488 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1949
timestamp 1626908933
transform 1 0 1488 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3213
timestamp 1626908933
transform 1 0 1488 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3916
timestamp 1626908933
transform 1 0 1488 0 1 5587
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1331
timestamp 1626908933
transform 1 0 1584 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1918
timestamp 1626908933
transform 1 0 1488 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3266
timestamp 1626908933
transform 1 0 1584 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3853
timestamp 1626908933
transform 1 0 1488 0 1 5587
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_684
timestamp 1626908933
transform 1 0 1440 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1406
timestamp 1626908933
transform 1 0 1440 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_579
timestamp 1626908933
transform 1 0 1056 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1177
timestamp 1626908933
transform 1 0 1056 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_528
timestamp 1626908933
transform 1 0 2208 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1519
timestamp 1626908933
transform 1 0 2208 0 -1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1921
timestamp 1626908933
transform 1 0 1968 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3856
timestamp 1626908933
transform 1 0 1968 0 1 5587
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_286
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_643
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_400
timestamp 1626908933
transform 1 0 2304 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1001
timestamp 1626908933
transform 1 0 2304 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1951
timestamp 1626908933
transform 1 0 2352 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3918
timestamp 1626908933
transform 1 0 2352 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3219
timestamp 1626908933
transform 1 0 2736 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1252
timestamp 1626908933
transform 1 0 2736 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_66
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_14
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_955
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_307
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_955
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_307
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3271
timestamp 1626908933
transform 1 0 2928 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1336
timestamp 1626908933
transform 1 0 2928 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3269
timestamp 1626908933
transform 1 0 3120 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3246
timestamp 1626908933
transform 1 0 3120 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1334
timestamp 1626908933
transform 1 0 3120 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1311
timestamp 1626908933
transform 1 0 3120 0 1 5439
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3218
timestamp 1626908933
transform 1 0 3120 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1251
timestamp 1626908933
transform 1 0 3120 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1711
timestamp 1626908933
transform 1 0 2976 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_720
timestamp 1626908933
transform 1 0 2976 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_319
timestamp 1626908933
transform 1 0 3216 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2286
timestamp 1626908933
transform 1 0 3216 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_1
timestamp 1626908933
transform 1 0 3072 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_4
timestamp 1626908933
transform 1 0 3072 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_631
timestamp 1626908933
transform 1 0 3552 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1353
timestamp 1626908933
transform 1 0 3552 0 -1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1221
timestamp 1626908933
transform 1 0 3984 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1230
timestamp 1626908933
transform 1 0 3888 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3188
timestamp 1626908933
transform 1 0 3984 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3197
timestamp 1626908933
transform 1 0 3888 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_345
timestamp 1626908933
transform 1 0 4080 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1293
timestamp 1626908933
transform 1 0 3888 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2280
timestamp 1626908933
transform 1 0 4080 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3228
timestamp 1626908933
transform 1 0 3888 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1151
timestamp 1626908933
transform 1 0 4272 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3118
timestamp 1626908933
transform 1 0 4272 0 1 5735
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1221
timestamp 1626908933
transform 1 0 4080 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3156
timestamp 1626908933
transform 1 0 4080 0 1 5735
box -29 -23 29 23
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_3
timestamp 1626908933
transform -1 0 4800 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_9
timestamp 1626908933
transform -1 0 4800 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_276
timestamp 1626908933
transform 1 0 4800 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_877
timestamp 1626908933
transform 1 0 4800 0 -1 6660
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1215
timestamp 1626908933
transform 1 0 4848 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1218
timestamp 1626908933
transform 1 0 4560 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3150
timestamp 1626908933
transform 1 0 4848 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3153
timestamp 1626908933
transform 1 0 4560 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_527
timestamp 1626908933
transform 1 0 4992 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1518
timestamp 1626908933
transform 1 0 4992 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1146
timestamp 1626908933
transform 1 0 4944 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3113
timestamp 1626908933
transform 1 0 4944 0 1 5883
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_283
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_931
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_283
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_931
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_609
timestamp 1626908933
transform 1 0 5088 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1331
timestamp 1626908933
transform 1 0 5088 0 -1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1154
timestamp 1626908933
transform 1 0 5808 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3121
timestamp 1626908933
transform 1 0 5808 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1225
timestamp 1626908933
transform 1 0 5808 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1409
timestamp 1626908933
transform 1 0 5808 0 1 5809
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3160
timestamp 1626908933
transform 1 0 5808 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3344
timestamp 1626908933
transform 1 0 5808 0 1 5809
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_52
timestamp 1626908933
transform -1 0 6240 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_114
timestamp 1626908933
transform -1 0 6240 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_484
timestamp 1626908933
transform 1 0 6432 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1082
timestamp 1626908933
transform 1 0 6432 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_275
timestamp 1626908933
transform 1 0 6240 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_876
timestamp 1626908933
transform 1 0 6240 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_125
timestamp 1626908933
transform 1 0 6384 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2092
timestamp 1626908933
transform 1 0 6384 0 1 5883
box -32 -32 32 32
use L1M1_PR  L1M1_PR_136
timestamp 1626908933
transform 1 0 6192 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2071
timestamp 1626908933
transform 1 0 6192 0 1 5883
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_98
timestamp 1626908933
transform 1 0 6816 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_29
timestamp 1626908933
transform 1 0 6816 0 -1 6660
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1327
timestamp 1626908933
transform 1 0 6672 0 1 5809
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3294
timestamp 1626908933
transform 1 0 6672 0 1 5809
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_401
timestamp 1626908933
transform 1 0 7296 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1002
timestamp 1626908933
transform 1 0 7296 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_285
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_642
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_721
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1712
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_259
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_907
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_259
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_907
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1743
timestamp 1626908933
transform 1 0 7920 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3710
timestamp 1626908933
transform 1 0 7920 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1527
timestamp 1626908933
transform 1 0 8208 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1939
timestamp 1626908933
transform 1 0 8208 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3494
timestamp 1626908933
transform 1 0 8208 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3906
timestamp 1626908933
transform 1 0 8208 0 1 5587
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1911
timestamp 1626908933
transform 1 0 8016 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3846
timestamp 1626908933
transform 1 0 8016 0 1 5587
box -29 -23 29 23
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_26
timestamp 1626908933
transform 1 0 7680 0 -1 6660
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_2
timestamp 1626908933
transform 1 0 7680 0 -1 6660
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_813
timestamp 1626908933
transform 1 0 8592 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2780
timestamp 1626908933
transform 1 0 8592 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_850
timestamp 1626908933
transform 1 0 8976 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2785
timestamp 1626908933
transform 1 0 8976 0 1 5439
box -29 -23 29 23
use M1M2_PR  M1M2_PR_27
timestamp 1626908933
transform 1 0 9264 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1994
timestamp 1626908933
transform 1 0 9264 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1614
timestamp 1626908933
transform 1 0 8304 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3549
timestamp 1626908933
transform 1 0 8304 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_28
timestamp 1626908933
transform 1 0 9264 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1963
timestamp 1626908933
transform 1 0 9264 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_402
timestamp 1626908933
transform 1 0 9984 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1003
timestamp 1626908933
transform 1 0 9984 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_722
timestamp 1626908933
transform 1 0 10176 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1713
timestamp 1626908933
transform 1 0 10176 0 -1 6660
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_235
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_883
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_235
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_883
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use M1M2_PR  M1M2_PR_911
timestamp 1626908933
transform 1 0 10416 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2878
timestamp 1626908933
transform 1 0 10416 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_963
timestamp 1626908933
transform 1 0 10320 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_969
timestamp 1626908933
transform 1 0 10416 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2898
timestamp 1626908933
transform 1 0 10320 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2904
timestamp 1626908933
transform 1 0 10416 0 1 5439
box -29 -23 29 23
use M1M2_PR  M1M2_PR_618
timestamp 1626908933
transform 1 0 10608 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_916
timestamp 1626908933
transform 1 0 10704 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2585
timestamp 1626908933
transform 1 0 10608 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2883
timestamp 1626908933
transform 1 0 10704 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_628
timestamp 1626908933
transform 1 0 10512 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2563
timestamp 1626908933
transform 1 0 10512 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_762
timestamp 1626908933
transform 1 0 10896 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2729
timestamp 1626908933
transform 1 0 10896 0 1 5513
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_29
timestamp 1626908933
transform 1 0 10272 0 -1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_4
timestamp 1626908933
transform 1 0 10272 0 -1 6660
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_149
timestamp 1626908933
transform 1 0 12048 0 1 5513
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2084
timestamp 1626908933
transform 1 0 12048 0 1 5513
box -29 -23 29 23
use M1M2_PR  M1M2_PR_131
timestamp 1626908933
transform 1 0 11568 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2098
timestamp 1626908933
transform 1 0 11568 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_143
timestamp 1626908933
transform 1 0 11568 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_631
timestamp 1626908933
transform 1 0 11760 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_793
timestamp 1626908933
transform 1 0 11664 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2078
timestamp 1626908933
transform 1 0 11568 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2566
timestamp 1626908933
transform 1 0 11760 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2728
timestamp 1626908933
transform 1 0 11664 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_630
timestamp 1626908933
transform 1 0 11952 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2597
timestamp 1626908933
transform 1 0 11952 0 1 5883
box -32 -32 32 32
use L1M1_PR  L1M1_PR_639
timestamp 1626908933
transform 1 0 11856 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2574
timestamp 1626908933
transform 1 0 11856 0 1 5883
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_211
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_859
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_211
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_859
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1517
timestamp 1626908933
transform 1 0 12576 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_526
timestamp 1626908933
transform 1 0 12576 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_641
timestamp 1626908933
transform 1 0 12480 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_284
timestamp 1626908933
transform 1 0 12480 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2101
timestamp 1626908933
transform 1 0 12720 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_134
timestamp 1626908933
transform 1 0 12720 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2587
timestamp 1626908933
transform 1 0 12912 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_620
timestamp 1626908933
transform 1 0 12912 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2564
timestamp 1626908933
transform 1 0 13008 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2558
timestamp 1626908933
transform 1 0 13104 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_629
timestamp 1626908933
transform 1 0 13008 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_623
timestamp 1626908933
transform 1 0 13104 0 1 5883
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2581
timestamp 1626908933
transform 1 0 13104 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_614
timestamp 1626908933
transform 1 0 13104 0 1 5883
box -32 -32 32 32
use L1M1_PR  L1M1_PR_146
timestamp 1626908933
transform 1 0 13296 0 1 5513
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2081
timestamp 1626908933
transform 1 0 13296 0 1 5513
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_464
timestamp 1626908933
transform 1 0 12672 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1186
timestamp 1626908933
transform 1 0 12672 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_32
timestamp 1626908933
transform 1 0 13440 0 -1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_7
timestamp 1626908933
transform 1 0 13440 0 -1 6660
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_2912
timestamp 1626908933
transform 1 0 14160 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2906
timestamp 1626908933
transform 1 0 14064 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_977
timestamp 1626908933
transform 1 0 14160 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_971
timestamp 1626908933
transform 1 0 14064 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2891
timestamp 1626908933
transform 1 0 14256 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2885
timestamp 1626908933
transform 1 0 13872 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_924
timestamp 1626908933
transform 1 0 14256 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_918
timestamp 1626908933
transform 1 0 13872 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_701
timestamp 1626908933
transform 1 0 15120 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2668
timestamp 1626908933
transform 1 0 15120 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_721
timestamp 1626908933
transform 1 0 15120 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2656
timestamp 1626908933
transform 1 0 15120 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_46
timestamp 1626908933
transform 1 0 15408 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1981
timestamp 1626908933
transform 1 0 15408 0 1 5587
box -29 -23 29 23
use M1M2_PR  M1M2_PR_612
timestamp 1626908933
transform 1 0 14736 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2579
timestamp 1626908933
transform 1 0 14736 0 1 5883
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_187
timestamp 1626908933
transform 1 0 14900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_835
timestamp 1626908933
transform 1 0 14900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_187
timestamp 1626908933
transform 1 0 14900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_835
timestamp 1626908933
transform 1 0 14900 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_620
timestamp 1626908933
transform 1 0 15312 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2555
timestamp 1626908933
transform 1 0 15312 0 1 5883
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_525
timestamp 1626908933
transform 1 0 15648 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1516
timestamp 1626908933
transform 1 0 15648 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_41
timestamp 1626908933
transform 1 0 15792 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_830
timestamp 1626908933
transform 1 0 15888 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2008
timestamp 1626908933
transform 1 0 15792 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2797
timestamp 1626908933
transform 1 0 15888 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_524
timestamp 1626908933
transform 1 0 16128 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1515
timestamp 1626908933
transform 1 0 16128 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1468
timestamp 1626908933
transform 1 0 16272 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3435
timestamp 1626908933
transform 1 0 16272 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1553
timestamp 1626908933
transform 1 0 16272 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3488
timestamp 1626908933
transform 1 0 16272 0 1 5439
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_394
timestamp 1626908933
transform 1 0 16224 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1116
timestamp 1626908933
transform 1 0 16224 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_307
timestamp 1626908933
transform 1 0 15744 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_905
timestamp 1626908933
transform 1 0 15744 0 -1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2809
timestamp 1626908933
transform 1 0 16464 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_874
timestamp 1626908933
transform 1 0 16464 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2802
timestamp 1626908933
transform 1 0 16368 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_835
timestamp 1626908933
transform 1 0 16368 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_523
timestamp 1626908933
transform 1 0 16992 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1514
timestamp 1626908933
transform 1 0 16992 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_44
timestamp 1626908933
transform 1 0 16752 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2011
timestamp 1626908933
transform 1 0 16752 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_50
timestamp 1626908933
transform 1 0 16752 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_869
timestamp 1626908933
transform 1 0 16656 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1985
timestamp 1626908933
transform 1 0 16752 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2804
timestamp 1626908933
transform 1 0 16656 0 1 5883
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_811
timestamp 1626908933
transform 1 0 17300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_163
timestamp 1626908933
transform 1 0 17300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_811
timestamp 1626908933
transform 1 0 17300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_163
timestamp 1626908933
transform 1 0 17300 0 1 5994
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3670
timestamp 1626908933
transform 1 0 17328 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1703
timestamp 1626908933
transform 1 0 17328 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_640
timestamp 1626908933
transform 1 0 17472 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_283
timestamp 1626908933
transform 1 0 17472 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_881
timestamp 1626908933
transform 1 0 17088 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_283
timestamp 1626908933
transform 1 0 17088 0 -1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_194
timestamp 1626908933
transform 1 0 17712 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2161
timestamp 1626908933
transform 1 0 17712 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_213
timestamp 1626908933
transform 1 0 17712 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2148
timestamp 1626908933
transform 1 0 17712 0 1 5439
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3665
timestamp 1626908933
transform 1 0 19056 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1698
timestamp 1626908933
transform 1 0 19056 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_47
timestamp 1626908933
transform -1 0 19872 0 -1 6660
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_23
timestamp 1626908933
transform -1 0 19872 0 -1 6660
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_1482
timestamp 1626908933
transform 1 0 19728 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1931
timestamp 1626908933
transform 1 0 19440 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3449
timestamp 1626908933
transform 1 0 19728 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3898
timestamp 1626908933
transform 1 0 19440 0 1 5587
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1569
timestamp 1626908933
transform 1 0 19824 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1898
timestamp 1626908933
transform 1 0 19536 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3504
timestamp 1626908933
transform 1 0 19824 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3833
timestamp 1626908933
transform 1 0 19536 0 1 5587
box -29 -23 29 23
use M1M2_PR  M1M2_PR_110
timestamp 1626908933
transform 1 0 20112 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2077
timestamp 1626908933
transform 1 0 20112 0 1 5883
box -32 -32 32 32
use L1M1_PR  L1M1_PR_124
timestamp 1626908933
transform 1 0 20112 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2059
timestamp 1626908933
transform 1 0 20112 0 1 5883
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_139
timestamp 1626908933
transform 1 0 19700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_787
timestamp 1626908933
transform 1 0 19700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_139
timestamp 1626908933
transform 1 0 19700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_787
timestamp 1626908933
transform 1 0 19700 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_223
timestamp 1626908933
transform 1 0 19872 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_821
timestamp 1626908933
transform 1 0 19872 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_50
timestamp 1626908933
transform -1 0 21024 0 -1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_11
timestamp 1626908933
transform -1 0 21024 0 -1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1004
timestamp 1626908933
transform 1 0 20256 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_403
timestamp 1626908933
transform 1 0 20256 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1010
timestamp 1626908933
transform 1 0 21024 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_288
timestamp 1626908933
transform 1 0 21024 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_2
timestamp 1626908933
transform 1 0 21792 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_71
timestamp 1626908933
transform 1 0 21792 0 -1 6660
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_763
timestamp 1626908933
transform 1 0 22100 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_115
timestamp 1626908933
transform 1 0 22100 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_763
timestamp 1626908933
transform 1 0 22100 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_115
timestamp 1626908933
transform 1 0 22100 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3830
timestamp 1626908933
transform 1 0 21936 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1895
timestamp 1626908933
transform 1 0 21936 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_282
timestamp 1626908933
transform 1 0 22464 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_639
timestamp 1626908933
transform 1 0 22464 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_404
timestamp 1626908933
transform 1 0 22272 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1005
timestamp 1626908933
transform 1 0 22272 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1437
timestamp 1626908933
transform 1 0 22320 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3404
timestamp 1626908933
transform 1 0 22320 0 1 5735
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1521
timestamp 1626908933
transform 1 0 22320 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3456
timestamp 1626908933
transform 1 0 22320 0 1 5735
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_522
timestamp 1626908933
transform 1 0 22560 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1513
timestamp 1626908933
transform 1 0 22560 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1442
timestamp 1626908933
transform 1 0 22800 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3409
timestamp 1626908933
transform 1 0 22800 0 1 5587
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1528
timestamp 1626908933
transform 1 0 22704 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3463
timestamp 1626908933
transform 1 0 22704 0 1 5587
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_175
timestamp 1626908933
transform 1 0 22656 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_773
timestamp 1626908933
transform 1 0 22656 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_10
timestamp 1626908933
transform -1 0 23616 0 -1 6660
box -38 -49 614 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_4
timestamp 1626908933
transform -1 0 23616 0 -1 6660
box -38 -49 614 715
use L1M1_PR  L1M1_PR_3829
timestamp 1626908933
transform 1 0 23088 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1894
timestamp 1626908933
transform 1 0 23088 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_28
timestamp 1626908933
transform 1 0 23616 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_5
timestamp 1626908933
transform 1 0 23616 0 -1 6660
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_739
timestamp 1626908933
transform 1 0 24500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_91
timestamp 1626908933
transform 1 0 24500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_739
timestamp 1626908933
transform 1 0 24500 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_91
timestamp 1626908933
transform 1 0 24500 0 1 5994
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2065
timestamp 1626908933
transform 1 0 24336 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_98
timestamp 1626908933
transform 1 0 24336 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_26
timestamp 1626908933
transform 1 0 24384 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_95
timestamp 1626908933
transform 1 0 24384 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_67
timestamp 1626908933
transform 1 0 24864 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_15
timestamp 1626908933
transform 1 0 24864 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_723
timestamp 1626908933
transform 1 0 25248 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1714
timestamp 1626908933
transform 1 0 25248 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1926
timestamp 1626908933
transform 1 0 25200 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3893
timestamp 1626908933
transform 1 0 25200 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_109
timestamp 1626908933
transform 1 0 24912 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2044
timestamp 1626908933
transform 1 0 24912 0 1 5883
box -29 -23 29 23
use M1M2_PR  M1M2_PR_726
timestamp 1626908933
transform 1 0 25392 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2693
timestamp 1626908933
transform 1 0 25392 0 1 5735
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_107
timestamp 1626908933
transform 1 0 25344 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_38
timestamp 1626908933
transform 1 0 25344 0 -1 6660
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2962
timestamp 1626908933
transform 1 0 26448 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2683
timestamp 1626908933
transform 1 0 26544 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1027
timestamp 1626908933
transform 1 0 26448 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_748
timestamp 1626908933
transform 1 0 26544 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2931
timestamp 1626908933
transform 1 0 26448 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_964
timestamp 1626908933
transform 1 0 26448 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_29
timestamp 1626908933
transform 1 0 25824 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_6
timestamp 1626908933
transform 1 0 25824 0 -1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_968
timestamp 1626908933
transform 1 0 26640 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1490
timestamp 1626908933
transform 1 0 26736 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2935
timestamp 1626908933
transform 1 0 26640 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3457
timestamp 1626908933
transform 1 0 26736 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1031
timestamp 1626908933
transform 1 0 26736 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1578
timestamp 1626908933
transform 1 0 26640 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2966
timestamp 1626908933
transform 1 0 26736 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3513
timestamp 1626908933
transform 1 0 26640 0 1 5439
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_724
timestamp 1626908933
transform 1 0 26592 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1715
timestamp 1626908933
transform 1 0 26592 0 -1 6660
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_715
timestamp 1626908933
transform 1 0 26900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_67
timestamp 1626908933
transform 1 0 26900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_715
timestamp 1626908933
transform 1 0 26900 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_67
timestamp 1626908933
transform 1 0 26900 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_91
timestamp 1626908933
transform 1 0 26688 0 -1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_29
timestamp 1626908933
transform 1 0 26688 0 -1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_725
timestamp 1626908933
transform 1 0 27360 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1716
timestamp 1626908933
transform 1 0 27360 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_92
timestamp 1626908933
transform 1 0 26976 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_690
timestamp 1626908933
transform 1 0 26976 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_875
timestamp 1626908933
transform 1 0 27552 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_274
timestamp 1626908933
transform 1 0 27552 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_638
timestamp 1626908933
transform 1 0 27456 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_281
timestamp 1626908933
transform 1 0 27456 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3648
timestamp 1626908933
transform 1 0 27696 0 1 5809
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1681
timestamp 1626908933
transform 1 0 27696 0 1 5809
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_855
timestamp 1626908933
transform 1 0 27744 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_133
timestamp 1626908933
transform 1 0 27744 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_521
timestamp 1626908933
transform 1 0 28896 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1512
timestamp 1626908933
transform 1 0 28896 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1782
timestamp 1626908933
transform 1 0 28752 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3749
timestamp 1626908933
transform 1 0 28752 0 1 5883
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_43
timestamp 1626908933
transform 1 0 29300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_691
timestamp 1626908933
transform 1 0 29300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_43
timestamp 1626908933
transform 1 0 29300 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_691
timestamp 1626908933
transform 1 0 29300 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_98
timestamp 1626908933
transform 1 0 28992 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_820
timestamp 1626908933
transform 1 0 28992 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_66
timestamp 1626908933
transform 1 0 28512 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_664
timestamp 1626908933
transform 1 0 28512 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_874
timestamp 1626908933
transform 1 0 29760 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_273
timestamp 1626908933
transform 1 0 29760 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_632
timestamp 1626908933
transform 1 0 29952 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_34
timestamp 1626908933
transform 1 0 29952 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_781
timestamp 1626908933
transform 1 0 30336 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_59
timestamp 1626908933
transform 1 0 30336 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_610
timestamp 1626908933
transform 1 0 31104 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_12
timestamp 1626908933
transform 1 0 31104 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_520
timestamp 1626908933
transform 1 0 31488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1511
timestamp 1626908933
transform 1 0 31488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_280
timestamp 1626908933
transform 1 0 31680 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_637
timestamp 1626908933
transform 1 0 31680 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_726
timestamp 1626908933
transform 1 0 31584 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1717
timestamp 1626908933
transform 1 0 31584 0 -1 6660
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_19
timestamp 1626908933
transform 1 0 31700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_667
timestamp 1626908933
transform 1 0 31700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_19
timestamp 1626908933
transform 1 0 31700 0 1 5994
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_667
timestamp 1626908933
transform 1 0 31700 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_405
timestamp 1626908933
transform 1 0 31776 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1006
timestamp 1626908933
transform 1 0 31776 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3747
timestamp 1626908933
transform 1 0 32016 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1780
timestamp 1626908933
transform 1 0 32016 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1718
timestamp 1626908933
transform 1 0 31968 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_727
timestamp 1626908933
transform 1 0 31968 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1719
timestamp 1626908933
transform 1 0 192 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_728
timestamp 1626908933
transform 1 0 192 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3917
timestamp 1626908933
transform 1 0 240 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1950
timestamp 1626908933
transform 1 0 240 0 1 6845
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_636
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_279
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1008
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1007
timestamp 1626908933
transform 1 0 0 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_407
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_406
timestamp 1626908933
transform 1 0 0 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_61
timestamp 1626908933
transform -1 0 960 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_123
timestamp 1626908933
transform -1 0 960 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_4
timestamp 1626908933
transform 1 0 960 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_9
timestamp 1626908933
transform 1 0 960 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_729
timestamp 1626908933
transform 1 0 1632 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1720
timestamp 1626908933
transform 1 0 1632 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1948
timestamp 1626908933
transform 1 0 1488 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3915
timestamp 1626908933
transform 1 0 1488 0 1 6845
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_643
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1291
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_643
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1291
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_578
timestamp 1626908933
transform 1 0 1248 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1176
timestamp 1626908933
transform 1 0 1248 0 1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_313
timestamp 1626908933
transform 1 0 1968 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2280
timestamp 1626908933
transform 1 0 1968 0 1 6401
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_272
timestamp 1626908933
transform 1 0 2400 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_873
timestamp 1626908933
transform 1 0 2400 0 1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_308
timestamp 1626908933
transform 1 0 2352 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1232
timestamp 1626908933
transform 1 0 2160 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2275
timestamp 1626908933
transform 1 0 2352 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3199
timestamp 1626908933
transform 1 0 2160 0 1 6771
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1315
timestamp 1626908933
transform 1 0 2160 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3250
timestamp 1626908933
transform 1 0 2160 0 1 6771
box -29 -23 29 23
use sky130_fd_sc_hs__a2bb2oi_1  sky130_fd_sc_hs__a2bb2oi_1_0
timestamp 1626908933
transform 1 0 1728 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__a2bb2oi_1  sky130_fd_sc_hs__a2bb2oi_1_1
timestamp 1626908933
transform 1 0 1728 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1510
timestamp 1626908933
transform 1 0 2592 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_519
timestamp 1626908933
transform 1 0 2592 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1379
timestamp 1626908933
transform 1 0 2688 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_657
timestamp 1626908933
transform 1 0 2688 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_332
timestamp 1626908933
transform 1 0 3024 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2267
timestamp 1626908933
transform 1 0 3024 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2272
timestamp 1626908933
transform 1 0 3216 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_337
timestamp 1626908933
transform 1 0 3216 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2285
timestamp 1626908933
transform 1 0 3312 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_318
timestamp 1626908933
transform 1 0 3312 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3229
timestamp 1626908933
transform 1 0 3408 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1294
timestamp 1626908933
transform 1 0 3408 0 1 6253
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3568
timestamp 1626908933
transform 1 0 3504 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1601
timestamp 1626908933
transform 1 0 3504 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1509
timestamp 1626908933
transform 1 0 3456 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_518
timestamp 1626908933
transform 1 0 3456 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_7
timestamp 1626908933
transform 1 0 3552 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_15
timestamp 1626908933
transform 1 0 3552 0 1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_1220
timestamp 1626908933
transform 1 0 3984 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3187
timestamp 1626908933
transform 1 0 3984 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1291
timestamp 1626908933
transform 1 0 4368 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1691
timestamp 1626908933
transform 1 0 4272 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3226
timestamp 1626908933
transform 1 0 4368 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3626
timestamp 1626908933
transform 1 0 4272 0 1 6549
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_619
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1267
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_619
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1267
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_623
timestamp 1626908933
transform 1 0 4224 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1345
timestamp 1626908933
transform 1 0 4224 0 1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_316
timestamp 1626908933
transform 1 0 4752 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1143
timestamp 1626908933
transform 1 0 4560 0 1 6475
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2283
timestamp 1626908933
transform 1 0 4752 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3110
timestamp 1626908933
transform 1 0 4560 0 1 6475
box -32 -32 32 32
use L1M1_PR  L1M1_PR_344
timestamp 1626908933
transform 1 0 4752 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1292
timestamp 1626908933
transform 1 0 4560 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2279
timestamp 1626908933
transform 1 0 4752 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3227
timestamp 1626908933
transform 1 0 4560 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3186
timestamp 1626908933
transform 1 0 4944 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3112
timestamp 1626908933
transform 1 0 4944 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1219
timestamp 1626908933
transform 1 0 4944 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1145
timestamp 1626908933
transform 1 0 4944 0 1 6327
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_635
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_278
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3111
timestamp 1626908933
transform 1 0 5040 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1144
timestamp 1626908933
transform 1 0 5040 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1009
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_408
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_57
timestamp 1626908933
transform 1 0 5280 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_119
timestamp 1626908933
transform 1 0 5280 0 1 6660
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2287
timestamp 1626908933
transform 1 0 5904 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_352
timestamp 1626908933
transform 1 0 5904 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2293
timestamp 1626908933
transform 1 0 5904 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_326
timestamp 1626908933
transform 1 0 5904 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3148
timestamp 1626908933
transform 1 0 6096 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1213
timestamp 1626908933
transform 1 0 6096 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2283
timestamp 1626908933
transform 1 0 6192 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_348
timestamp 1626908933
transform 1 0 6192 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2289
timestamp 1626908933
transform 1 0 6192 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_322
timestamp 1626908933
transform 1 0 6192 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3146
timestamp 1626908933
transform 1 0 6000 0 1 6475
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1211
timestamp 1626908933
transform 1 0 6000 0 1 6475
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1214
timestamp 1626908933
transform 1 0 5616 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3149
timestamp 1626908933
transform 1 0 5616 0 1 6771
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_124
timestamp 1626908933
transform 1 0 5952 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_55
timestamp 1626908933
transform 1 0 5952 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_16
timestamp 1626908933
transform 1 0 5568 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_68
timestamp 1626908933
transform 1 0 5568 0 1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_124
timestamp 1626908933
transform 1 0 6384 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2091
timestamp 1626908933
transform 1 0 6384 0 1 6327
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_595
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1243
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_595
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1243
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_135
timestamp 1626908933
transform 1 0 6864 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_808
timestamp 1626908933
transform 1 0 7152 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2070
timestamp 1626908933
transform 1 0 6864 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2743
timestamp 1626908933
transform 1 0 7152 0 1 6549
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_38
timestamp 1626908933
transform -1 0 7488 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_100
timestamp 1626908933
transform -1 0 7488 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_579
timestamp 1626908933
transform 1 0 6432 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1301
timestamp 1626908933
transform 1 0 6432 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_517
timestamp 1626908933
transform 1 0 7488 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1508
timestamp 1626908933
transform 1 0 7488 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_776
timestamp 1626908933
transform 1 0 7248 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_777
timestamp 1626908933
transform 1 0 7248 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2743
timestamp 1626908933
transform 1 0 7248 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2744
timestamp 1626908933
transform 1 0 7248 0 1 6549
box -32 -32 32 32
use L1M1_PR  L1M1_PR_807
timestamp 1626908933
transform 1 0 7536 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2742
timestamp 1626908933
transform 1 0 7536 0 1 6771
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_516
timestamp 1626908933
transform 1 0 7968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1507
timestamp 1626908933
transform 1 0 7968 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1742
timestamp 1626908933
transform 1 0 7920 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3709
timestamp 1626908933
transform 1 0 7920 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1564
timestamp 1626908933
transform 1 0 7728 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3499
timestamp 1626908933
transform 1 0 7728 0 1 6401
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_472
timestamp 1626908933
transform 1 0 7584 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1070
timestamp 1626908933
transform 1 0 7584 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_26
timestamp 1626908933
transform 1 0 8064 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_88
timestamp 1626908933
transform 1 0 8064 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3845
timestamp 1626908933
transform 1 0 8112 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1910
timestamp 1626908933
transform 1 0 8112 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3908
timestamp 1626908933
transform 1 0 8112 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3493
timestamp 1626908933
transform 1 0 8208 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1941
timestamp 1626908933
transform 1 0 8112 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1526
timestamp 1626908933
transform 1 0 8208 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_271
timestamp 1626908933
transform 1 0 8448 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_872
timestamp 1626908933
transform 1 0 8448 0 1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1735
timestamp 1626908933
transform 1 0 8400 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3702
timestamp 1626908933
transform 1 0 8400 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1613
timestamp 1626908933
transform 1 0 8304 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3548
timestamp 1626908933
transform 1 0 8304 0 1 6771
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1476
timestamp 1626908933
transform 1 0 8688 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3443
timestamp 1626908933
transform 1 0 8688 0 1 6401
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_571
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1219
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_571
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1219
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_449
timestamp 1626908933
transform 1 0 8640 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1047
timestamp 1626908933
transform 1 0 8640 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_71
timestamp 1626908933
transform -1 0 9312 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_9
timestamp 1626908933
transform -1 0 9312 0 1 6660
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1993
timestamp 1626908933
transform 1 0 9264 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_26
timestamp 1626908933
transform 1 0 9264 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1506
timestamp 1626908933
transform 1 0 9312 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_515
timestamp 1626908933
transform 1 0 9312 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1035
timestamp 1626908933
transform 1 0 9408 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_437
timestamp 1626908933
transform 1 0 9408 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1961
timestamp 1626908933
transform 1 0 9936 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_26
timestamp 1626908933
transform 1 0 9936 0 1 6105
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1721
timestamp 1626908933
transform 1 0 9888 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1505
timestamp 1626908933
transform 1 0 9792 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_730
timestamp 1626908933
transform 1 0 9888 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_514
timestamp 1626908933
transform 1 0 9792 0 1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3545
timestamp 1626908933
transform 1 0 10320 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1610
timestamp 1626908933
transform 1 0 10320 0 1 6253
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1010
timestamp 1626908933
transform 1 0 10080 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_409
timestamp 1626908933
transform 1 0 10080 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_634
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_277
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_14
timestamp 1626908933
transform 1 0 10272 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_83
timestamp 1626908933
transform 1 0 10272 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_410
timestamp 1626908933
transform 1 0 10752 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1011
timestamp 1626908933
transform 1 0 10752 0 1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_617
timestamp 1626908933
transform 1 0 10608 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2584
timestamp 1626908933
transform 1 0 10608 0 1 6845
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1906
timestamp 1626908933
transform 1 0 10608 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3841
timestamp 1626908933
transform 1 0 10608 0 1 6401
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_731
timestamp 1626908933
transform 1 0 10944 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1722
timestamp 1626908933
transform 1 0 10944 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_0
timestamp 1626908933
transform 1 0 11040 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_2
timestamp 1626908933
transform 1 0 11040 0 1 6660
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1522
timestamp 1626908933
transform 1 0 11088 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3489
timestamp 1626908933
transform 1 0 11088 0 1 6253
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_547
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1195
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_547
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1195
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_411
timestamp 1626908933
transform 1 0 11520 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1012
timestamp 1626908933
transform 1 0 11520 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_732
timestamp 1626908933
transform 1 0 11712 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1723
timestamp 1626908933
transform 1 0 11712 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_130
timestamp 1626908933
transform 1 0 11568 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2097
timestamp 1626908933
transform 1 0 11568 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_99
timestamp 1626908933
transform 1 0 11808 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_30
timestamp 1626908933
transform 1 0 11808 0 1 6660
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2561
timestamp 1626908933
transform 1 0 11952 0 1 6845
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2076
timestamp 1626908933
transform 1 0 12432 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_626
timestamp 1626908933
transform 1 0 11952 0 1 6845
box -29 -23 29 23
use L1M1_PR  L1M1_PR_141
timestamp 1626908933
transform 1 0 12432 0 1 6105
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_871
timestamp 1626908933
transform 1 0 12288 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_270
timestamp 1626908933
transform 1 0 12288 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_970
timestamp 1626908933
transform 1 0 12480 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_372
timestamp 1626908933
transform 1 0 12480 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_8
timestamp 1626908933
transform 1 0 12864 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_0
timestamp 1626908933
transform 1 0 12864 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3539
timestamp 1626908933
transform 1 0 13392 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1604
timestamp 1626908933
transform 1 0 13392 0 1 6549
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2583
timestamp 1626908933
transform 1 0 13008 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_616
timestamp 1626908933
transform 1 0 13008 0 1 6845
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1169
timestamp 1626908933
transform 1 0 13248 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_447
timestamp 1626908933
transform 1 0 13248 0 1 6660
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1171
timestamp 1626908933
transform 1 0 13700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_523
timestamp 1626908933
transform 1 0 13700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1171
timestamp 1626908933
transform 1 0 13700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_523
timestamp 1626908933
transform 1 0 13700 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3840
timestamp 1626908933
transform 1 0 13776 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1905
timestamp 1626908933
transform 1 0 13776 0 1 6401
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_269
timestamp 1626908933
transform 1 0 14400 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_870
timestamp 1626908933
transform 1 0 14400 0 1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1517
timestamp 1626908933
transform 1 0 14544 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1936
timestamp 1626908933
transform 1 0 14544 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3484
timestamp 1626908933
transform 1 0 14544 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3903
timestamp 1626908933
transform 1 0 14544 0 1 6401
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_336
timestamp 1626908933
transform 1 0 14592 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_934
timestamp 1626908933
transform 1 0 14592 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_4
timestamp 1626908933
transform 1 0 14016 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_12
timestamp 1626908933
transform 1 0 14016 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_276
timestamp 1626908933
transform 1 0 14976 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_633
timestamp 1626908933
transform 1 0 14976 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_268
timestamp 1626908933
transform 1 0 15072 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_869
timestamp 1626908933
transform 1 0 15072 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_513
timestamp 1626908933
transform 1 0 15264 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1504
timestamp 1626908933
transform 1 0 15264 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_142
timestamp 1626908933
transform 1 0 15408 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2109
timestamp 1626908933
transform 1 0 15408 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_414
timestamp 1626908933
transform 1 0 15360 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1136
timestamp 1626908933
transform 1 0 15360 0 1 6660
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1147
timestamp 1626908933
transform 1 0 16100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_499
timestamp 1626908933
transform 1 0 16100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1147
timestamp 1626908933
transform 1 0 16100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_499
timestamp 1626908933
transform 1 0 16100 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2091
timestamp 1626908933
transform 1 0 15600 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_156
timestamp 1626908933
transform 1 0 15600 0 1 6549
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_80
timestamp 1626908933
transform 1 0 16128 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_19
timestamp 1626908933
transform 1 0 16128 0 1 6660
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2810
timestamp 1626908933
transform 1 0 16368 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_875
timestamp 1626908933
transform 1 0 16368 0 1 6771
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2801
timestamp 1626908933
transform 1 0 16368 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_834
timestamp 1626908933
transform 1 0 16368 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_868
timestamp 1626908933
transform 1 0 16416 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_267
timestamp 1626908933
transform 1 0 16416 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_26
timestamp 1626908933
transform 1 0 17376 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_1
timestamp 1626908933
transform 1 0 17376 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1107
timestamp 1626908933
transform 1 0 16608 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_385
timestamp 1626908933
transform 1 0 16608 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2063
timestamp 1626908933
transform 1 0 17616 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_128
timestamp 1626908933
transform 1 0 17616 0 1 6549
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2084
timestamp 1626908933
transform 1 0 17712 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_117
timestamp 1626908933
transform 1 0 17712 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1503
timestamp 1626908933
transform 1 0 17856 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_512
timestamp 1626908933
transform 1 0 17856 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1083
timestamp 1626908933
transform 1 0 17952 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_361
timestamp 1626908933
transform 1 0 17952 0 1 6660
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1123
timestamp 1626908933
transform 1 0 18500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_475
timestamp 1626908933
transform 1 0 18500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1123
timestamp 1626908933
transform 1 0 18500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_475
timestamp 1626908933
transform 1 0 18500 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_8
timestamp 1626908933
transform 1 0 18720 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_0
timestamp 1626908933
transform 1 0 18720 0 1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_3664
timestamp 1626908933
transform 1 0 19056 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1697
timestamp 1626908933
transform 1 0 19056 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3455
timestamp 1626908933
transform 1 0 19344 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1520
timestamp 1626908933
transform 1 0 19344 0 1 6771
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2768
timestamp 1626908933
transform 1 0 19152 0 1 6179
box -32 -32 32 32
use M1M2_PR  M1M2_PR_801
timestamp 1626908933
transform 1 0 19152 0 1 6179
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3834
timestamp 1626908933
transform 1 0 19440 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1899
timestamp 1626908933
transform 1 0 19440 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3897
timestamp 1626908933
transform 1 0 19440 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1930
timestamp 1626908933
transform 1 0 19440 0 1 6327
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1502
timestamp 1626908933
transform 1 0 19392 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_511
timestamp 1626908933
transform 1 0 19392 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3402
timestamp 1626908933
transform 1 0 19728 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3401
timestamp 1626908933
transform 1 0 19728 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1435
timestamp 1626908933
transform 1 0 19728 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1434
timestamp 1626908933
transform 1 0 19728 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_275
timestamp 1626908933
transform 1 0 19968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_632
timestamp 1626908933
transform 1 0 19968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_510
timestamp 1626908933
transform 1 0 19872 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1501
timestamp 1626908933
transform 1 0 19872 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_109
timestamp 1626908933
transform 1 0 20112 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2076
timestamp 1626908933
transform 1 0 20112 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1519
timestamp 1626908933
transform 1 0 19824 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3454
timestamp 1626908933
transform 1 0 19824 0 1 6401
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_309
timestamp 1626908933
transform 1 0 20064 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1031
timestamp 1626908933
transform 1 0 20064 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_230
timestamp 1626908933
transform 1 0 19488 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_828
timestamp 1626908933
transform 1 0 19488 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_121
timestamp 1626908933
transform 1 0 20496 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_942
timestamp 1626908933
transform 1 0 20592 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2056
timestamp 1626908933
transform 1 0 20496 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2877
timestamp 1626908933
transform 1 0 20592 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2768
timestamp 1626908933
transform 1 0 20784 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_833
timestamp 1626908933
transform 1 0 20784 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2859
timestamp 1626908933
transform 1 0 20688 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_892
timestamp 1626908933
transform 1 0 20688 0 1 6401
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1099
timestamp 1626908933
transform 1 0 20900 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_451
timestamp 1626908933
transform 1 0 20900 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1099
timestamp 1626908933
transform 1 0 20900 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_451
timestamp 1626908933
transform 1 0 20900 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3457
timestamp 1626908933
transform 1 0 20976 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1522
timestamp 1626908933
transform 1 0 20976 0 1 6105
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1500
timestamp 1626908933
transform 1 0 20832 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_509
timestamp 1626908933
transform 1 0 20832 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_205
timestamp 1626908933
transform 1 0 20928 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_803
timestamp 1626908933
transform 1 0 20928 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2508
timestamp 1626908933
transform 1 0 21840 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_573
timestamp 1626908933
transform 1 0 21840 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2536
timestamp 1626908933
transform 1 0 21072 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2504
timestamp 1626908933
transform 1 0 21840 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_569
timestamp 1626908933
transform 1 0 21072 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_537
timestamp 1626908933
transform 1 0 21840 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1009
timestamp 1626908933
transform 1 0 21312 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_287
timestamp 1626908933
transform 1 0 21312 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2473
timestamp 1626908933
transform 1 0 21936 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_538
timestamp 1626908933
transform 1 0 21936 0 1 6549
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1499
timestamp 1626908933
transform 1 0 22080 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_508
timestamp 1626908933
transform 1 0 22080 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_65
timestamp 1626908933
transform -1 0 23328 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_3
timestamp 1626908933
transform -1 0 23328 0 1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3403
timestamp 1626908933
transform 1 0 22320 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2505
timestamp 1626908933
transform 1 0 22320 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1436
timestamp 1626908933
transform 1 0 22320 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_538
timestamp 1626908933
transform 1 0 22320 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_979
timestamp 1626908933
transform 1 0 22176 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_257
timestamp 1626908933
transform 1 0 22176 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2475
timestamp 1626908933
transform 1 0 23088 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_540
timestamp 1626908933
transform 1 0 23088 0 1 6549
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2542
timestamp 1626908933
transform 1 0 23088 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_575
timestamp 1626908933
transform 1 0 23088 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_572
timestamp 1626908933
transform 1 0 23280 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_580
timestamp 1626908933
transform 1 0 23184 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2507
timestamp 1626908933
transform 1 0 23280 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2515
timestamp 1626908933
transform 1 0 23184 0 1 6401
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_427
timestamp 1626908933
transform 1 0 23300 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1075
timestamp 1626908933
transform 1 0 23300 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_427
timestamp 1626908933
transform 1 0 23300 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1075
timestamp 1626908933
transform 1 0 23300 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_507
timestamp 1626908933
transform 1 0 23328 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1498
timestamp 1626908933
transform 1 0 23328 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_791
timestamp 1626908933
transform 1 0 23760 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2758
timestamp 1626908933
transform 1 0 23760 0 1 6105
box -32 -32 32 32
use L1M1_PR  L1M1_PR_198
timestamp 1626908933
transform 1 0 23664 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_825
timestamp 1626908933
transform 1 0 23472 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2133
timestamp 1626908933
transform 1 0 23664 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2760
timestamp 1626908933
transform 1 0 23472 0 1 6105
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_225
timestamp 1626908933
transform 1 0 23424 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_947
timestamp 1626908933
transform 1 0 23424 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_111
timestamp 1626908933
transform 1 0 24144 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2046
timestamp 1626908933
transform 1 0 24144 0 1 6771
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_4
timestamp 1626908933
transform 1 0 24192 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_66
timestamp 1626908933
transform 1 0 24192 0 1 6660
box -38 -49 326 715
use M1M2_PR  M1M2_PR_97
timestamp 1626908933
transform 1 0 24432 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2064
timestamp 1626908933
transform 1 0 24432 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_110
timestamp 1626908933
transform 1 0 24432 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_823
timestamp 1626908933
transform 1 0 24528 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2045
timestamp 1626908933
transform 1 0 24432 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2758
timestamp 1626908933
transform 1 0 24528 0 1 6105
box -29 -23 29 23
use M1M2_PR  M1M2_PR_96
timestamp 1626908933
transform 1 0 24432 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2063
timestamp 1626908933
transform 1 0 24432 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_506
timestamp 1626908933
transform 1 0 24480 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1497
timestamp 1626908933
transform 1 0 24480 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_137
timestamp 1626908933
transform 1 0 24576 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_735
timestamp 1626908933
transform 1 0 24576 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_274
timestamp 1626908933
transform 1 0 24960 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_631
timestamp 1626908933
transform 1 0 24960 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_125
timestamp 1626908933
transform 1 0 25056 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_723
timestamp 1626908933
transform 1 0 25056 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_197
timestamp 1626908933
transform 1 0 25296 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2132
timestamp 1626908933
transform 1 0 25296 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_725
timestamp 1626908933
transform 1 0 25392 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2692
timestamp 1626908933
transform 1 0 25392 0 1 6549
box -32 -32 32 32
use L1M1_PR  L1M1_PR_749
timestamp 1626908933
transform 1 0 25488 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2684
timestamp 1626908933
transform 1 0 25488 0 1 6549
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_403
timestamp 1626908933
transform 1 0 25700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1051
timestamp 1626908933
transform 1 0 25700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_403
timestamp 1626908933
transform 1 0 25700 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1051
timestamp 1626908933
transform 1 0 25700 0 1 6660
box -100 -49 100 49
use M1M2_PR  M1M2_PR_180
timestamp 1626908933
transform 1 0 26256 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2147
timestamp 1626908933
transform 1 0 26256 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_963
timestamp 1626908933
transform 1 0 26448 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2930
timestamp 1626908933
transform 1 0 26448 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_967
timestamp 1626908933
transform 1 0 26640 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2934
timestamp 1626908933
transform 1 0 26640 0 1 6105
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1025
timestamp 1626908933
transform 1 0 26928 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1030
timestamp 1626908933
transform 1 0 26832 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2960
timestamp 1626908933
transform 1 0 26928 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2965
timestamp 1626908933
transform 1 0 26832 0 1 6105
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_505
timestamp 1626908933
transform 1 0 27648 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1496
timestamp 1626908933
transform 1 0 27648 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_44
timestamp 1626908933
transform 1 0 25440 0 1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_19
timestamp 1626908933
transform 1 0 25440 0 1 6660
box -38 -49 2246 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1027
timestamp 1626908933
transform 1 0 28100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_379
timestamp 1626908933
transform 1 0 28100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1027
timestamp 1626908933
transform 1 0 28100 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_379
timestamp 1626908933
transform 1 0 28100 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_854
timestamp 1626908933
transform 1 0 27744 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_132
timestamp 1626908933
transform 1 0 27744 0 1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3752
timestamp 1626908933
transform 1 0 29136 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1785
timestamp 1626908933
transform 1 0 29136 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1495
timestamp 1626908933
transform 1 0 28896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_504
timestamp 1626908933
transform 1 0 28896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_663
timestamp 1626908933
transform 1 0 28512 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_65
timestamp 1626908933
transform 1 0 28512 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_819
timestamp 1626908933
transform 1 0 28992 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_97
timestamp 1626908933
transform 1 0 28992 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_867
timestamp 1626908933
transform 1 0 29760 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_866
timestamp 1626908933
transform 1 0 30048 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_266
timestamp 1626908933
transform 1 0 29760 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_265
timestamp 1626908933
transform 1 0 30048 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_630
timestamp 1626908933
transform 1 0 29952 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_273
timestamp 1626908933
transform 1 0 29952 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1494
timestamp 1626908933
transform 1 0 30240 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_503
timestamp 1626908933
transform 1 0 30240 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_780
timestamp 1626908933
transform 1 0 30336 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_58
timestamp 1626908933
transform 1 0 30336 0 1 6660
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1003
timestamp 1626908933
transform 1 0 30500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_355
timestamp 1626908933
transform 1 0 30500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1003
timestamp 1626908933
transform 1 0 30500 0 1 6660
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_355
timestamp 1626908933
transform 1 0 30500 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1493
timestamp 1626908933
transform 1 0 31104 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_502
timestamp 1626908933
transform 1 0 31104 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_740
timestamp 1626908933
transform 1 0 31200 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_18
timestamp 1626908933
transform 1 0 31200 0 1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3750
timestamp 1626908933
transform 1 0 31920 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1783
timestamp 1626908933
transform 1 0 31920 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1724
timestamp 1626908933
transform 1 0 31968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_733
timestamp 1626908933
transform 1 0 31968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_264
timestamp 1626908933
transform 1 0 0 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_865
timestamp 1626908933
transform 1 0 0 0 -1 7992
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3280
timestamp 1626908933
transform 1 0 624 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1345
timestamp 1626908933
transform 1 0 624 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3227
timestamp 1626908933
transform 1 0 720 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1260
timestamp 1626908933
transform 1 0 720 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2277
timestamp 1626908933
transform 1 0 816 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_342
timestamp 1626908933
transform 1 0 816 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3279
timestamp 1626908933
transform 1 0 624 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1344
timestamp 1626908933
transform 1 0 624 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3226
timestamp 1626908933
transform 1 0 720 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1259
timestamp 1626908933
transform 1 0 720 0 1 7215
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_978
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_330
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_978
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_330
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_716
timestamp 1626908933
transform 1 0 192 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1438
timestamp 1626908933
transform 1 0 192 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1263
timestamp 1626908933
transform 1 0 1104 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3230
timestamp 1626908933
transform 1 0 1104 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_341
timestamp 1626908933
transform 1 0 1008 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1348
timestamp 1626908933
transform 1 0 1104 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1919
timestamp 1626908933
transform 1 0 912 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2276
timestamp 1626908933
transform 1 0 1008 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3283
timestamp 1626908933
transform 1 0 1104 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3854
timestamp 1626908933
transform 1 0 912 0 1 6919
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_57
timestamp 1626908933
transform 1 0 1344 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_118
timestamp 1626908933
transform 1 0 1344 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_501
timestamp 1626908933
transform 1 0 1632 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1492
timestamp 1626908933
transform 1 0 1632 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1335
timestamp 1626908933
transform 1 0 1488 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3270
timestamp 1626908933
transform 1 0 1488 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_577
timestamp 1626908933
transform 1 0 960 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1175
timestamp 1626908933
transform 1 0 960 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_315
timestamp 1626908933
transform 1 0 1872 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1244
timestamp 1626908933
transform 1 0 1776 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2282
timestamp 1626908933
transform 1 0 1872 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3211
timestamp 1626908933
transform 1 0 1776 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_340
timestamp 1626908933
transform 1 0 1872 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1326
timestamp 1626908933
transform 1 0 1776 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2275
timestamp 1626908933
transform 1 0 1872 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3261
timestamp 1626908933
transform 1 0 1776 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3852
timestamp 1626908933
transform 1 0 2256 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1917
timestamp 1626908933
transform 1 0 2256 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3737
timestamp 1626908933
transform 1 0 2160 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1770
timestamp 1626908933
transform 1 0 2160 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2269
timestamp 1626908933
transform 1 0 2448 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_334
timestamp 1626908933
transform 1 0 2448 0 1 7067
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2274
timestamp 1626908933
transform 1 0 2352 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_307
timestamp 1626908933
transform 1 0 2352 0 1 7067
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_629
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_272
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_662
timestamp 1626908933
transform 1 0 1728 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1384
timestamp 1626908933
transform 1 0 1728 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1013
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_412
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_954
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_306
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_954
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_306
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1725
timestamp 1626908933
transform 1 0 2784 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_734
timestamp 1626908933
transform 1 0 2784 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3217
timestamp 1626908933
transform 1 0 3120 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1250
timestamp 1626908933
transform 1 0 3120 0 1 7437
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_864
timestamp 1626908933
transform 1 0 3168 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_263
timestamp 1626908933
transform 1 0 3168 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_116
timestamp 1626908933
transform 1 0 2880 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_55
timestamp 1626908933
transform 1 0 2880 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_648
timestamp 1626908933
transform 1 0 3360 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1370
timestamp 1626908933
transform 1 0 3360 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_331
timestamp 1626908933
transform 1 0 3696 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2298
timestamp 1626908933
transform 1 0 3696 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_356
timestamp 1626908933
transform 1 0 3888 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1210
timestamp 1626908933
transform 1 0 3888 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1784
timestamp 1626908933
transform 1 0 3984 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2291
timestamp 1626908933
transform 1 0 3888 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3145
timestamp 1626908933
transform 1 0 3888 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3719
timestamp 1626908933
transform 1 0 3984 0 1 7215
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_262
timestamp 1626908933
transform 1 0 4128 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_863
timestamp 1626908933
transform 1 0 4128 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_735
timestamp 1626908933
transform 1 0 4320 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1726
timestamp 1626908933
transform 1 0 4320 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1140
timestamp 1626908933
transform 1 0 4080 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1141
timestamp 1626908933
transform 1 0 4080 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3107
timestamp 1626908933
transform 1 0 4080 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3108
timestamp 1626908933
transform 1 0 4080 0 1 7067
box -32 -32 32 32
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_6
timestamp 1626908933
transform -1 0 4800 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_14
timestamp 1626908933
transform -1 0 4800 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_500
timestamp 1626908933
transform 1 0 4800 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1491
timestamp 1626908933
transform 1 0 4800 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1208
timestamp 1626908933
transform 1 0 4464 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3143
timestamp 1626908933
transform 1 0 4464 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1217
timestamp 1626908933
transform 1 0 5136 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1218
timestamp 1626908933
transform 1 0 4944 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3184
timestamp 1626908933
transform 1 0 5136 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3185
timestamp 1626908933
transform 1 0 4944 0 1 6993
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_282
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_930
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_282
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_930
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_608
timestamp 1626908933
transform 1 0 5280 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1330
timestamp 1626908933
transform 1 0 5280 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_511
timestamp 1626908933
transform 1 0 4896 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1109
timestamp 1626908933
transform 1 0 4896 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3225
timestamp 1626908933
transform 1 0 5328 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3224
timestamp 1626908933
transform 1 0 5424 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1290
timestamp 1626908933
transform 1 0 5328 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1289
timestamp 1626908933
transform 1 0 5424 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3115
timestamp 1626908933
transform 1 0 5520 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1148
timestamp 1626908933
transform 1 0 5520 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_325
timestamp 1626908933
transform 1 0 5904 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2292
timestamp 1626908933
transform 1 0 5904 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_261
timestamp 1626908933
transform 1 0 6048 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_862
timestamp 1626908933
transform 1 0 6048 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_499
timestamp 1626908933
transform 1 0 6240 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1490
timestamp 1626908933
transform 1 0 6240 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_351
timestamp 1626908933
transform 1 0 6000 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1216
timestamp 1626908933
transform 1 0 6096 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2286
timestamp 1626908933
transform 1 0 6000 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3151
timestamp 1626908933
transform 1 0 6096 0 1 7215
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_578
timestamp 1626908933
transform 1 0 6336 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1300
timestamp 1626908933
transform 1 0 6336 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2876
timestamp 1626908933
transform 1 0 7056 0 1 7141
box -32 -32 32 32
use M1M2_PR  M1M2_PR_909
timestamp 1626908933
transform 1 0 7056 0 1 7141
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_95
timestamp 1626908933
transform 1 0 7104 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_34
timestamp 1626908933
transform 1 0 7104 0 -1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2895
timestamp 1626908933
transform 1 0 7344 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2892
timestamp 1626908933
transform 1 0 7248 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_960
timestamp 1626908933
transform 1 0 7344 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_957
timestamp 1626908933
transform 1 0 7248 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2873
timestamp 1626908933
transform 1 0 7344 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_906
timestamp 1626908933
transform 1 0 7344 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1727
timestamp 1626908933
transform 1 0 7392 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_736
timestamp 1626908933
transform 1 0 7392 0 -1 7992
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_906
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_258
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_906
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_258
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_628
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_271
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_861
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_260
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_498
timestamp 1626908933
transform 1 0 7776 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1489
timestamp 1626908933
transform 1 0 7776 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_559
timestamp 1626908933
transform 1 0 7872 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1281
timestamp 1626908933
transform 1 0 7872 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2889
timestamp 1626908933
transform 1 0 8112 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2741
timestamp 1626908933
transform 1 0 8208 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_954
timestamp 1626908933
transform 1 0 8112 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_806
timestamp 1626908933
transform 1 0 8208 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2742
timestamp 1626908933
transform 1 0 8208 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_775
timestamp 1626908933
transform 1 0 8208 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2894
timestamp 1626908933
transform 1 0 8496 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2739
timestamp 1626908933
transform 1 0 9072 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_959
timestamp 1626908933
transform 1 0 8496 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_804
timestamp 1626908933
transform 1 0 9072 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1046
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_448
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1261
timestamp 1626908933
transform 1 0 9024 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_539
timestamp 1626908933
transform 1 0 9024 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1962
timestamp 1626908933
transform 1 0 9264 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_27
timestamp 1626908933
transform 1 0 9264 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1992
timestamp 1626908933
transform 1 0 9264 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_25
timestamp 1626908933
transform 1 0 9264 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2093
timestamp 1626908933
transform 1 0 9744 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_126
timestamp 1626908933
transform 1 0 9744 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2577
timestamp 1626908933
transform 1 0 9168 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_642
timestamp 1626908933
transform 1 0 9168 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2601
timestamp 1626908933
transform 1 0 9456 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_634
timestamp 1626908933
transform 1 0 9456 0 1 7215
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_12
timestamp 1626908933
transform -1 0 10176 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_74
timestamp 1626908933
transform -1 0 10176 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_28
timestamp 1626908933
transform 1 0 10032 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1995
timestamp 1626908933
transform 1 0 10032 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_137
timestamp 1626908933
transform 1 0 10320 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2072
timestamp 1626908933
transform 1 0 10320 0 1 6993
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_234
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_882
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_234
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_882
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2587
timestamp 1626908933
transform 1 0 10416 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_652
timestamp 1626908933
transform 1 0 10416 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2609
timestamp 1626908933
transform 1 0 10416 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_642
timestamp 1626908933
transform 1 0 10416 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2586
timestamp 1626908933
transform 1 0 10416 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_651
timestamp 1626908933
transform 1 0 10416 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2608
timestamp 1626908933
transform 1 0 10416 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_641
timestamp 1626908933
transform 1 0 10416 0 1 7437
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1014
timestamp 1626908933
transform 1 0 10560 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_413
timestamp 1626908933
transform 1 0 10560 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_62
timestamp 1626908933
transform 1 0 10752 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_1
timestamp 1626908933
transform 1 0 10752 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_17
timestamp 1626908933
transform 1 0 10176 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_69
timestamp 1626908933
transform 1 0 10176 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_860
timestamp 1626908933
transform 1 0 11040 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_259
timestamp 1626908933
transform 1 0 11040 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_497
timestamp 1626908933
transform 1 0 11232 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1488
timestamp 1626908933
transform 1 0 11232 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_30
timestamp 1626908933
transform 1 0 11280 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1965
timestamp 1626908933
transform 1 0 11280 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_129
timestamp 1626908933
transform 1 0 11568 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2096
timestamp 1626908933
transform 1 0 11568 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_636
timestamp 1626908933
transform 1 0 11472 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2571
timestamp 1626908933
transform 1 0 11472 0 1 7215
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_399
timestamp 1626908933
transform 1 0 11328 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_997
timestamp 1626908933
transform 1 0 11328 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_5
timestamp 1626908933
transform 1 0 11712 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_67
timestamp 1626908933
transform 1 0 11712 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_35
timestamp 1626908933
transform 1 0 12336 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_627
timestamp 1626908933
transform 1 0 11760 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2002
timestamp 1626908933
transform 1 0 12336 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2594
timestamp 1626908933
transform 1 0 11760 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_142
timestamp 1626908933
transform 1 0 11856 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2077
timestamp 1626908933
transform 1 0 11856 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_629
timestamp 1626908933
transform 1 0 11952 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2596
timestamp 1626908933
transform 1 0 11952 0 1 7437
box -32 -32 32 32
use L1M1_PR  L1M1_PR_638
timestamp 1626908933
transform 1 0 12144 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2573
timestamp 1626908933
transform 1 0 12144 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_18
timestamp 1626908933
transform 1 0 12096 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_70
timestamp 1626908933
transform 1 0 12096 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_270
timestamp 1626908933
transform 1 0 12480 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_627
timestamp 1626908933
transform 1 0 12480 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_414
timestamp 1626908933
transform 1 0 12576 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1015
timestamp 1626908933
transform 1 0 12576 0 -1 7992
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_210
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_858
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_210
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_858
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use L1M1_PR  L1M1_PR_36
timestamp 1626908933
transform 1 0 12912 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_764
timestamp 1626908933
transform 1 0 13008 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1971
timestamp 1626908933
transform 1 0 12912 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2699
timestamp 1626908933
transform 1 0 13008 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_8
timestamp 1626908933
transform 1 0 12768 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_70
timestamp 1626908933
transform 1 0 12768 0 -1 7992
box -38 -49 326 715
use M1M2_PR  M1M2_PR_613
timestamp 1626908933
transform 1 0 13104 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2580
timestamp 1626908933
transform 1 0 13104 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_622
timestamp 1626908933
transform 1 0 13104 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2557
timestamp 1626908933
transform 1 0 13104 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_624
timestamp 1626908933
transform 1 0 13200 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2559
timestamp 1626908933
transform 1 0 13200 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_741
timestamp 1626908933
transform 1 0 13296 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2708
timestamp 1626908933
transform 1 0 13296 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_618
timestamp 1626908933
transform 1 0 13200 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2553
timestamp 1626908933
transform 1 0 13200 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2707
timestamp 1626908933
transform 1 0 13296 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_740
timestamp 1626908933
transform 1 0 13296 0 1 7437
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1487
timestamp 1626908933
transform 1 0 13056 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_496
timestamp 1626908933
transform 1 0 13056 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_495
timestamp 1626908933
transform 1 0 13536 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1486
timestamp 1626908933
transform 1 0 13536 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_354
timestamp 1626908933
transform 1 0 13152 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_952
timestamp 1626908933
transform 1 0 13152 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_1
timestamp 1626908933
transform 1 0 13632 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_5
timestamp 1626908933
transform 1 0 13632 0 -1 7992
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2550
timestamp 1626908933
transform 1 0 13776 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_615
timestamp 1626908933
transform 1 0 13776 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2576
timestamp 1626908933
transform 1 0 13776 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_609
timestamp 1626908933
transform 1 0 13776 0 1 7215
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_494
timestamp 1626908933
transform 1 0 14208 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1485
timestamp 1626908933
transform 1 0 14208 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_605
timestamp 1626908933
transform 1 0 14064 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_606
timestamp 1626908933
transform 1 0 14064 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2572
timestamp 1626908933
transform 1 0 14064 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2573
timestamp 1626908933
transform 1 0 14064 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_614
timestamp 1626908933
transform 1 0 14064 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2549
timestamp 1626908933
transform 1 0 14064 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2698
timestamp 1626908933
transform 1 0 14256 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_763
timestamp 1626908933
transform 1 0 14256 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2652
timestamp 1626908933
transform 1 0 14352 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_717
timestamp 1626908933
transform 1 0 14352 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2665
timestamp 1626908933
transform 1 0 14352 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_698
timestamp 1626908933
transform 1 0 14352 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2546
timestamp 1626908933
transform 1 0 14448 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_611
timestamp 1626908933
transform 1 0 14448 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3483
timestamp 1626908933
transform 1 0 14544 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1516
timestamp 1626908933
transform 1 0 14544 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2890
timestamp 1626908933
transform 1 0 14256 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_923
timestamp 1626908933
transform 1 0 14256 0 1 7585
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_432
timestamp 1626908933
transform 1 0 14304 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1154
timestamp 1626908933
transform 1 0 14304 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_141
timestamp 1626908933
transform 1 0 15408 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_604
timestamp 1626908933
transform 1 0 15216 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2108
timestamp 1626908933
transform 1 0 15408 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2571
timestamp 1626908933
transform 1 0 15216 0 1 7215
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_834
timestamp 1626908933
transform 1 0 14900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_186
timestamp 1626908933
transform 1 0 14900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_834
timestamp 1626908933
transform 1 0 14900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_186
timestamp 1626908933
transform 1 0 14900 0 1 7326
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2570
timestamp 1626908933
transform 1 0 15216 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_603
timestamp 1626908933
transform 1 0 15216 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2889
timestamp 1626908933
transform 1 0 14928 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_922
timestamp 1626908933
transform 1 0 14928 0 1 7585
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3538
timestamp 1626908933
transform 1 0 15120 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1603
timestamp 1626908933
transform 1 0 15120 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2909
timestamp 1626908933
transform 1 0 15504 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_974
timestamp 1626908933
transform 1 0 15504 0 1 7585
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_15
timestamp 1626908933
transform 1 0 15072 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_54
timestamp 1626908933
transform 1 0 15072 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_493
timestamp 1626908933
transform 1 0 15648 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1484
timestamp 1626908933
transform 1 0 15648 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_829
timestamp 1626908933
transform 1 0 15888 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2796
timestamp 1626908933
transform 1 0 15888 0 1 6919
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_492
timestamp 1626908933
transform 1 0 16128 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1483
timestamp 1626908933
transform 1 0 16128 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_610
timestamp 1626908933
transform 1 0 16272 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_870
timestamp 1626908933
transform 1 0 16176 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2545
timestamp 1626908933
transform 1 0 16272 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2805
timestamp 1626908933
transform 1 0 16176 0 1 6919
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_306
timestamp 1626908933
transform 1 0 15744 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_904
timestamp 1626908933
transform 1 0 15744 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_2
timestamp 1626908933
transform -1 0 16704 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_27
timestamp 1626908933
transform -1 0 16704 0 -1 7992
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1987
timestamp 1626908933
transform 1 0 16368 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_52
timestamp 1626908933
transform 1 0 16368 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_47
timestamp 1626908933
transform 1 0 16656 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2014
timestamp 1626908933
transform 1 0 16656 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_153
timestamp 1626908933
transform 1 0 17328 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2088
timestamp 1626908933
transform 1 0 17328 0 1 6993
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_162
timestamp 1626908933
transform 1 0 17300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_810
timestamp 1626908933
transform 1 0 17300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_162
timestamp 1626908933
transform 1 0 17300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_810
timestamp 1626908933
transform 1 0 17300 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_384
timestamp 1626908933
transform 1 0 16704 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1106
timestamp 1626908933
transform 1 0 16704 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1482
timestamp 1626908933
transform 1 0 17568 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_491
timestamp 1626908933
transform 1 0 17568 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_626
timestamp 1626908933
transform 1 0 17472 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_269
timestamp 1626908933
transform 1 0 17472 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1983
timestamp 1626908933
transform 1 0 17616 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_48
timestamp 1626908933
transform 1 0 17616 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2569
timestamp 1626908933
transform 1 0 17616 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2083
timestamp 1626908933
transform 1 0 17712 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_602
timestamp 1626908933
transform 1 0 17616 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_116
timestamp 1626908933
transform 1 0 17712 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2529
timestamp 1626908933
transform 1 0 17808 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_594
timestamp 1626908933
transform 1 0 17808 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2554
timestamp 1626908933
transform 1 0 17808 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_587
timestamp 1626908933
transform 1 0 17808 0 1 7215
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_490
timestamp 1626908933
transform 1 0 18048 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1481
timestamp 1626908933
transform 1 0 18048 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_360
timestamp 1626908933
transform 1 0 18144 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1082
timestamp 1626908933
transform 1 0 18144 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_272
timestamp 1626908933
transform 1 0 17664 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_870
timestamp 1626908933
transform 1 0 17664 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2770
timestamp 1626908933
transform 1 0 19056 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2062
timestamp 1626908933
transform 1 0 19056 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_835
timestamp 1626908933
transform 1 0 19056 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_127
timestamp 1626908933
transform 1 0 19056 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1480
timestamp 1626908933
transform 1 0 18912 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_489
timestamp 1626908933
transform 1 0 18912 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_840
timestamp 1626908933
transform 1 0 19008 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_242
timestamp 1626908933
transform 1 0 19008 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2767
timestamp 1626908933
transform 1 0 19152 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2766
timestamp 1626908933
transform 1 0 19152 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_800
timestamp 1626908933
transform 1 0 19152 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_799
timestamp 1626908933
transform 1 0 19152 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_115
timestamp 1626908933
transform 1 0 19536 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2082
timestamp 1626908933
transform 1 0 19536 0 1 6993
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_138
timestamp 1626908933
transform 1 0 19700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_786
timestamp 1626908933
transform 1 0 19700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_138
timestamp 1626908933
transform 1 0 19700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_786
timestamp 1626908933
transform 1 0 19700 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_488
timestamp 1626908933
transform 1 0 20160 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1479
timestamp 1626908933
transform 1 0 20160 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_331
timestamp 1626908933
transform 1 0 19392 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1053
timestamp 1626908933
transform 1 0 19392 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2769
timestamp 1626908933
transform 1 0 20400 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_834
timestamp 1626908933
transform 1 0 20400 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1478
timestamp 1626908933
transform 1 0 20544 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_487
timestamp 1626908933
transform 1 0 20544 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1024
timestamp 1626908933
transform 1 0 20640 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_302
timestamp 1626908933
transform 1 0 20640 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_72
timestamp 1626908933
transform -1 0 20544 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_11
timestamp 1626908933
transform -1 0 20544 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_6
timestamp 1626908933
transform 1 0 21408 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_0
timestamp 1626908933
transform 1 0 21408 0 -1 7992
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_762
timestamp 1626908933
transform 1 0 22100 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_114
timestamp 1626908933
transform 1 0 22100 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_762
timestamp 1626908933
transform 1 0 22100 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_114
timestamp 1626908933
transform 1 0 22100 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1477
timestamp 1626908933
transform 1 0 21984 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_486
timestamp 1626908933
transform 1 0 21984 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_784
timestamp 1626908933
transform 1 0 22080 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_186
timestamp 1626908933
transform 1 0 22080 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2502
timestamp 1626908933
transform 1 0 22800 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_535
timestamp 1626908933
transform 1 0 22800 0 1 7215
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_978
timestamp 1626908933
transform 1 0 22560 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_256
timestamp 1626908933
transform 1 0 22560 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_625
timestamp 1626908933
transform 1 0 22464 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_268
timestamp 1626908933
transform 1 0 22464 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_577
timestamp 1626908933
transform 1 0 22992 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2544
timestamp 1626908933
transform 1 0 22992 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_583
timestamp 1626908933
transform 1 0 22992 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2518
timestamp 1626908933
transform 1 0 22992 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_574
timestamp 1626908933
transform 1 0 23088 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2541
timestamp 1626908933
transform 1 0 23088 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_579
timestamp 1626908933
transform 1 0 23280 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2514
timestamp 1626908933
transform 1 0 23280 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_577
timestamp 1626908933
transform 1 0 23184 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2512
timestamp 1626908933
transform 1 0 23184 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_536
timestamp 1626908933
transform 1 0 22992 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2471
timestamp 1626908933
transform 1 0 22992 0 1 7215
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_859
timestamp 1626908933
transform 1 0 23328 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_258
timestamp 1626908933
transform 1 0 23328 0 -1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_572
timestamp 1626908933
transform 1 0 23472 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2539
timestamp 1626908933
transform 1 0 23472 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_162
timestamp 1626908933
transform 1 0 23520 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_760
timestamp 1626908933
transform 1 0 23520 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_575
timestamp 1626908933
transform 1 0 24336 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_750
timestamp 1626908933
transform 1 0 24432 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2510
timestamp 1626908933
transform 1 0 24336 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2685
timestamp 1626908933
transform 1 0 24432 0 1 6993
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_90
timestamp 1626908933
transform 1 0 24500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_738
timestamp 1626908933
transform 1 0 24500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_90
timestamp 1626908933
transform 1 0 24500 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_738
timestamp 1626908933
transform 1 0 24500 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_224
timestamp 1626908933
transform 1 0 23904 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_946
timestamp 1626908933
transform 1 0 23904 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1476
timestamp 1626908933
transform 1 0 24672 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_485
timestamp 1626908933
transform 1 0 24672 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_734
timestamp 1626908933
transform 1 0 24768 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_136
timestamp 1626908933
transform 1 0 24768 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_724
timestamp 1626908933
transform 1 0 25392 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1493
timestamp 1626908933
transform 1 0 25488 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1925
timestamp 1626908933
transform 1 0 25200 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2691
timestamp 1626908933
transform 1 0 25392 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3460
timestamp 1626908933
transform 1 0 25488 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3892
timestamp 1626908933
transform 1 0 25200 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1579
timestamp 1626908933
transform 1 0 25488 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3514
timestamp 1626908933
transform 1 0 25488 0 1 7067
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_191
timestamp 1626908933
transform 1 0 25152 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_913
timestamp 1626908933
transform 1 0 25152 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3828
timestamp 1626908933
transform 1 0 25776 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1893
timestamp 1626908933
transform 1 0 25776 0 1 6919
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_858
timestamp 1626908933
transform 1 0 25920 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_257
timestamp 1626908933
transform 1 0 25920 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_707
timestamp 1626908933
transform 1 0 26112 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_109
timestamp 1626908933
transform 1 0 26112 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_886
timestamp 1626908933
transform 1 0 26496 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_164
timestamp 1626908933
transform 1 0 26496 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_179
timestamp 1626908933
transform 1 0 26736 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2146
timestamp 1626908933
transform 1 0 26736 0 1 7215
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_66
timestamp 1626908933
transform 1 0 26900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_714
timestamp 1626908933
transform 1 0 26900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_66
timestamp 1626908933
transform 1 0 26900 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_714
timestamp 1626908933
transform 1 0 26900 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_484
timestamp 1626908933
transform 1 0 27264 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_737
timestamp 1626908933
transform 1 0 27360 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1475
timestamp 1626908933
transform 1 0 27264 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1728
timestamp 1626908933
transform 1 0 27360 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2128
timestamp 1626908933
transform 1 0 27600 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_193
timestamp 1626908933
transform 1 0 27600 0 1 7215
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_857
timestamp 1626908933
transform 1 0 27552 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_256
timestamp 1626908933
transform 1 0 27552 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_624
timestamp 1626908933
transform 1 0 27456 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_267
timestamp 1626908933
transform 1 0 27456 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3647
timestamp 1626908933
transform 1 0 27696 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1680
timestamp 1626908933
transform 1 0 27696 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_853
timestamp 1626908933
transform 1 0 27744 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_131
timestamp 1626908933
transform 1 0 27744 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_483
timestamp 1626908933
transform 1 0 28896 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1474
timestamp 1626908933
transform 1 0 28896 0 -1 7992
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_42
timestamp 1626908933
transform 1 0 29300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_690
timestamp 1626908933
transform 1 0 29300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_42
timestamp 1626908933
transform 1 0 29300 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_690
timestamp 1626908933
transform 1 0 29300 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_96
timestamp 1626908933
transform 1 0 28992 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_818
timestamp 1626908933
transform 1 0 28992 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_64
timestamp 1626908933
transform 1 0 28512 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_662
timestamp 1626908933
transform 1 0 28512 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_856
timestamp 1626908933
transform 1 0 29760 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_255
timestamp 1626908933
transform 1 0 29760 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_631
timestamp 1626908933
transform 1 0 29952 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_33
timestamp 1626908933
transform 1 0 29952 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_779
timestamp 1626908933
transform 1 0 30336 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_57
timestamp 1626908933
transform 1 0 30336 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_609
timestamp 1626908933
transform 1 0 31104 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_11
timestamp 1626908933
transform 1 0 31104 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_482
timestamp 1626908933
transform 1 0 31488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1473
timestamp 1626908933
transform 1 0 31488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_266
timestamp 1626908933
transform 1 0 31680 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_623
timestamp 1626908933
transform 1 0 31680 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_738
timestamp 1626908933
transform 1 0 31584 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1729
timestamp 1626908933
transform 1 0 31584 0 -1 7992
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_18
timestamp 1626908933
transform 1 0 31700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_666
timestamp 1626908933
transform 1 0 31700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_18
timestamp 1626908933
transform 1 0 31700 0 1 7326
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_666
timestamp 1626908933
transform 1 0 31700 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_415
timestamp 1626908933
transform 1 0 31776 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1016
timestamp 1626908933
transform 1 0 31776 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1730
timestamp 1626908933
transform 1 0 31968 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_739
timestamp 1626908933
transform 1 0 31968 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_265
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_622
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_254
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_416
timestamp 1626908933
transform 1 0 0 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_855
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1017
timestamp 1626908933
transform 1 0 0 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_740
timestamp 1626908933
transform 1 0 192 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1731
timestamp 1626908933
transform 1 0 192 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_481
timestamp 1626908933
transform 1 0 576 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1472
timestamp 1626908933
transform 1 0 576 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1258
timestamp 1626908933
transform 1 0 720 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3225
timestamp 1626908933
transform 1 0 720 0 1 7733
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_696
timestamp 1626908933
transform 1 0 672 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1418
timestamp 1626908933
transform 1 0 672 0 1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1262
timestamp 1626908933
transform 1 0 1104 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3229
timestamp 1626908933
transform 1 0 1104 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_58
timestamp 1626908933
transform -1 0 1728 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_119
timestamp 1626908933
transform -1 0 1728 0 1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_1343
timestamp 1626908933
transform 1 0 1392 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1347
timestamp 1626908933
transform 1 0 1488 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3278
timestamp 1626908933
transform 1 0 1392 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3282
timestamp 1626908933
transform 1 0 1488 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1227
timestamp 1626908933
transform 1 0 1680 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1228
timestamp 1626908933
transform 1 0 1584 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3162
timestamp 1626908933
transform 1 0 1680 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3163
timestamp 1626908933
transform 1 0 1584 0 1 8177
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_642
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1290
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_642
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1290
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use M1M2_PR  M1M2_PR_314
timestamp 1626908933
transform 1 0 1872 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1156
timestamp 1626908933
transform 1 0 1872 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1157
timestamp 1626908933
transform 1 0 1872 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2281
timestamp 1626908933
transform 1 0 1872 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3123
timestamp 1626908933
transform 1 0 1872 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3124
timestamp 1626908933
transform 1 0 1872 0 1 7881
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_60
timestamp 1626908933
transform 1 0 2112 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_122
timestamp 1626908933
transform 1 0 2112 0 1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3722
timestamp 1626908933
transform 1 0 2352 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3720
timestamp 1626908933
transform 1 0 2160 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3161
timestamp 1626908933
transform 1 0 2448 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1787
timestamp 1626908933
transform 1 0 2352 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1785
timestamp 1626908933
transform 1 0 2160 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1226
timestamp 1626908933
transform 1 0 2448 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3736
timestamp 1626908933
transform 1 0 2160 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1769
timestamp 1626908933
transform 1 0 2160 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_121
timestamp 1626908933
transform 1 0 2400 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_60
timestamp 1626908933
transform 1 0 2400 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_19
timestamp 1626908933
transform 1 0 1728 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_71
timestamp 1626908933
transform 1 0 1728 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_480
timestamp 1626908933
transform 1 0 2688 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1471
timestamp 1626908933
transform 1 0 2688 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1158
timestamp 1626908933
transform 1 0 2640 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1159
timestamp 1626908933
transform 1 0 2640 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3125
timestamp 1626908933
transform 1 0 2640 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3126
timestamp 1626908933
transform 1 0 2640 0 1 7881
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1231
timestamp 1626908933
transform 1 0 2640 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3166
timestamp 1626908933
transform 1 0 2640 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1772
timestamp 1626908933
transform 1 0 2736 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3739
timestamp 1626908933
transform 1 0 2736 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_479
timestamp 1626908933
transform 1 0 3168 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1470
timestamp 1626908933
transform 1 0 3168 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_338
timestamp 1626908933
transform 1 0 2928 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1229
timestamp 1626908933
transform 1 0 3120 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1333
timestamp 1626908933
transform 1 0 3120 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2273
timestamp 1626908933
transform 1 0 2928 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3164
timestamp 1626908933
transform 1 0 3120 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3268
timestamp 1626908933
transform 1 0 3120 0 1 7733
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3216
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3215
timestamp 1626908933
transform 1 0 3312 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1249
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1248
timestamp 1626908933
transform 1 0 3312 0 1 8103
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1732
timestamp 1626908933
transform 1 0 3264 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_741
timestamp 1626908933
transform 1 0 3264 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3267
timestamp 1626908933
transform 1 0 3504 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2266
timestamp 1626908933
transform 1 0 3408 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1332
timestamp 1626908933
transform 1 0 3504 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_331
timestamp 1626908933
transform 1 0 3408 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_6
timestamp 1626908933
transform 1 0 3360 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_1
timestamp 1626908933
transform 1 0 3360 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_547
timestamp 1626908933
transform 1 0 2784 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1145
timestamp 1626908933
transform 1 0 2784 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_253
timestamp 1626908933
transform 1 0 3648 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_854
timestamp 1626908933
transform 1 0 3648 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1149
timestamp 1626908933
transform 1 0 4368 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1150
timestamp 1626908933
transform 1 0 4272 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3116
timestamp 1626908933
transform 1 0 4368 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3117
timestamp 1626908933
transform 1 0 4272 0 1 7659
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_618
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1266
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_618
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1266
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_527
timestamp 1626908933
transform 1 0 3840 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1125
timestamp 1626908933
transform 1 0 3840 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_3
timestamp 1626908933
transform 1 0 4224 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_11
timestamp 1626908933
transform 1 0 4224 0 1 7992
box -38 -49 710 715
use L1M1_PR  L1M1_PR_3155
timestamp 1626908933
transform 1 0 4464 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3152
timestamp 1626908933
transform 1 0 4560 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1220
timestamp 1626908933
transform 1 0 4464 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1217
timestamp 1626908933
transform 1 0 4560 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2361
timestamp 1626908933
transform 1 0 4752 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_426
timestamp 1626908933
transform 1 0 4752 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3154
timestamp 1626908933
transform 1 0 4464 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2362
timestamp 1626908933
transform 1 0 4560 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1219
timestamp 1626908933
transform 1 0 4464 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_427
timestamp 1626908933
transform 1 0 4560 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2398
timestamp 1626908933
transform 1 0 4944 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2397
timestamp 1626908933
transform 1 0 4944 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_431
timestamp 1626908933
transform 1 0 4944 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_430
timestamp 1626908933
transform 1 0 4944 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1733
timestamp 1626908933
transform 1 0 4896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_742
timestamp 1626908933
transform 1 0 4896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_621
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_264
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3183
timestamp 1626908933
transform 1 0 5136 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1216
timestamp 1626908933
transform 1 0 5136 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_853
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_252
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_607
timestamp 1626908933
transform 1 0 5280 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1329
timestamp 1626908933
transform 1 0 5280 0 1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3114
timestamp 1626908933
transform 1 0 5520 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2396
timestamp 1626908933
transform 1 0 5520 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1147
timestamp 1626908933
transform 1 0 5520 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_429
timestamp 1626908933
transform 1 0 5520 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_49
timestamp 1626908933
transform 1 0 6336 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_24
timestamp 1626908933
transform 1 0 6336 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1734
timestamp 1626908933
transform 1 0 6240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_743
timestamp 1626908933
transform 1 0 6240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_852
timestamp 1626908933
transform 1 0 6048 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_251
timestamp 1626908933
transform 1 0 6048 0 1 7992
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1242
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_594
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1242
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_594
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3223
timestamp 1626908933
transform 1 0 6384 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1288
timestamp 1626908933
transform 1 0 6384 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3296
timestamp 1626908933
transform 1 0 6480 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1329
timestamp 1626908933
transform 1 0 6480 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3343
timestamp 1626908933
transform 1 0 6576 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1408
timestamp 1626908933
transform 1 0 6576 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2090
timestamp 1626908933
transform 1 0 6864 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2087
timestamp 1626908933
transform 1 0 6960 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_123
timestamp 1626908933
transform 1 0 6864 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_120
timestamp 1626908933
transform 1 0 6960 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1469
timestamp 1626908933
transform 1 0 6816 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_478
timestamp 1626908933
transform 1 0 6816 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2872
timestamp 1626908933
transform 1 0 7056 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_905
timestamp 1626908933
transform 1 0 7056 0 1 7733
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2886
timestamp 1626908933
transform 1 0 7152 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_951
timestamp 1626908933
transform 1 0 7152 0 1 7733
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_567
timestamp 1626908933
transform 1 0 6912 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1289
timestamp 1626908933
transform 1 0 6912 0 1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_908
timestamp 1626908933
transform 1 0 7248 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2875
timestamp 1626908933
transform 1 0 7248 0 1 7881
box -32 -32 32 32
use L1M1_PR  L1M1_PR_132
timestamp 1626908933
transform 1 0 7344 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_955
timestamp 1626908933
transform 1 0 7344 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2067
timestamp 1626908933
transform 1 0 7344 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2890
timestamp 1626908933
transform 1 0 7344 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_131
timestamp 1626908933
transform 1 0 7728 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2066
timestamp 1626908933
transform 1 0 7728 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_82
timestamp 1626908933
transform 1 0 7680 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_13
timestamp 1626908933
transform 1 0 7680 0 1 7992
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2733
timestamp 1626908933
transform 1 0 8112 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_798
timestamp 1626908933
transform 1 0 8112 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2741
timestamp 1626908933
transform 1 0 8208 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_774
timestamp 1626908933
transform 1 0 8208 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1052
timestamp 1626908933
transform 1 0 8160 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_454
timestamp 1626908933
transform 1 0 8160 0 1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_798
timestamp 1626908933
transform 1 0 8688 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2765
timestamp 1626908933
transform 1 0 8688 0 1 7733
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_570
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1218
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_570
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1218
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2767
timestamp 1626908933
transform 1 0 8592 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_832
timestamp 1626908933
transform 1 0 8592 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2764
timestamp 1626908933
transform 1 0 8688 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_797
timestamp 1626908933
transform 1 0 8688 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2740
timestamp 1626908933
transform 1 0 8784 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2732
timestamp 1626908933
transform 1 0 8880 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_805
timestamp 1626908933
transform 1 0 8784 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_797
timestamp 1626908933
transform 1 0 8880 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1959
timestamp 1626908933
transform 1 0 9072 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_24
timestamp 1626908933
transform 1 0 9072 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1990
timestamp 1626908933
transform 1 0 9072 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_23
timestamp 1626908933
transform 1 0 9072 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_14
timestamp 1626908933
transform -1 0 9216 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_29
timestamp 1626908933
transform -1 0 9216 0 1 7992
box -38 -49 710 715
use M1M2_PR  M1M2_PR_24
timestamp 1626908933
transform 1 0 9264 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1991
timestamp 1626908933
transform 1 0 9264 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_29
timestamp 1626908933
transform 1 0 9168 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1964
timestamp 1626908933
transform 1 0 9168 0 1 8103
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_263
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_620
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_29
timestamp 1626908933
transform 1 0 9936 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1996
timestamp 1626908933
transform 1 0 9936 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_647
timestamp 1626908933
transform 1 0 9936 0 1 7807
box -29 -23 29 23
use L1M1_PR  L1M1_PR_831
timestamp 1626908933
transform 1 0 9840 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2582
timestamp 1626908933
transform 1 0 9936 0 1 7807
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2766
timestamp 1626908933
transform 1 0 9840 0 1 7733
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_526
timestamp 1626908933
transform 1 0 9216 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1248
timestamp 1626908933
transform 1 0 9216 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1967
timestamp 1626908933
transform 1 0 10032 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_32
timestamp 1626908933
transform 1 0 10032 0 1 7659
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1024
timestamp 1626908933
transform 1 0 10080 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_426
timestamp 1626908933
transform 1 0 10080 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1242
timestamp 1626908933
transform 1 0 10464 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_520
timestamp 1626908933
transform 1 0 10464 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2579
timestamp 1626908933
transform 1 0 10992 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1966
timestamp 1626908933
transform 1 0 10992 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_644
timestamp 1626908933
transform 1 0 10992 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_31
timestamp 1626908933
transform 1 0 10992 0 1 7733
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2603
timestamp 1626908933
transform 1 0 10992 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_636
timestamp 1626908933
transform 1 0 10992 0 1 7881
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_477
timestamp 1626908933
transform 1 0 11232 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1468
timestamp 1626908933
transform 1 0 11232 0 1 7992
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_546
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1194
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_546
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1194
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use M1M2_PR  M1M2_PR_626
timestamp 1626908933
transform 1 0 11760 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_638
timestamp 1626908933
transform 1 0 11664 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2593
timestamp 1626908933
transform 1 0 11760 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2605
timestamp 1626908933
transform 1 0 11664 0 1 7807
box -32 -32 32 32
use L1M1_PR  L1M1_PR_632
timestamp 1626908933
transform 1 0 11856 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_635
timestamp 1626908933
transform 1 0 11760 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2567
timestamp 1626908933
transform 1 0 11856 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2570
timestamp 1626908933
transform 1 0 11760 0 1 7733
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_487
timestamp 1626908933
transform 1 0 11712 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1209
timestamp 1626908933
transform 1 0 11712 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_398
timestamp 1626908933
transform 1 0 11328 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_996
timestamp 1626908933
transform 1 0 11328 0 1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_623
timestamp 1626908933
transform 1 0 11952 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_628
timestamp 1626908933
transform 1 0 12144 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2590
timestamp 1626908933
transform 1 0 11952 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2595
timestamp 1626908933
transform 1 0 12144 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_613
timestamp 1626908933
transform 1 0 11952 0 1 7807
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2548
timestamp 1626908933
transform 1 0 11952 0 1 7807
box -29 -23 29 23
use M1M2_PR  M1M2_PR_34
timestamp 1626908933
transform 1 0 12336 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2001
timestamp 1626908933
transform 1 0 12336 0 1 7659
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_250
timestamp 1626908933
transform 1 0 12480 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_851
timestamp 1626908933
transform 1 0 12480 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_476
timestamp 1626908933
transform 1 0 12672 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1467
timestamp 1626908933
transform 1 0 12672 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1972
timestamp 1626908933
transform 1 0 12816 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_37
timestamp 1626908933
transform 1 0 12816 0 1 7659
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1735
timestamp 1626908933
transform 1 0 12768 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_744
timestamp 1626908933
transform 1 0 12768 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2572
timestamp 1626908933
transform 1 0 13008 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2560
timestamp 1626908933
transform 1 0 13008 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_637
timestamp 1626908933
transform 1 0 13008 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_625
timestamp 1626908933
transform 1 0 13008 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2592
timestamp 1626908933
transform 1 0 13008 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2582
timestamp 1626908933
transform 1 0 13008 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_625
timestamp 1626908933
transform 1 0 13008 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_615
timestamp 1626908933
transform 1 0 13008 0 1 7659
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_249
timestamp 1626908933
transform 1 0 13440 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_850
timestamp 1626908933
transform 1 0 13440 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_665
timestamp 1626908933
transform 1 0 13392 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2632
timestamp 1626908933
transform 1 0 13392 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_680
timestamp 1626908933
transform 1 0 13392 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2615
timestamp 1626908933
transform 1 0 13392 0 1 8251
box -29 -23 29 23
use sky130_fd_sc_hs__nor4_1  sky130_fd_sc_hs__nor4_1_0
timestamp 1626908933
transform -1 0 13440 0 1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__nor4_1  sky130_fd_sc_hs__nor4_1_2
timestamp 1626908933
transform -1 0 13440 0 1 7992
box -38 -49 614 715
use M1M2_PR  M1M2_PR_608
timestamp 1626908933
transform 1 0 13776 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2575
timestamp 1626908933
transform 1 0 13776 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_612
timestamp 1626908933
transform 1 0 13680 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2547
timestamp 1626908933
transform 1 0 13680 0 1 7733
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_522
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1170
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_522
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1170
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_446
timestamp 1626908933
transform 1 0 13632 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1168
timestamp 1626908933
transform 1 0 13632 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_605
timestamp 1626908933
transform 1 0 14160 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_617
timestamp 1626908933
transform 1 0 14064 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_621
timestamp 1626908933
transform 1 0 14160 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2540
timestamp 1626908933
transform 1 0 14160 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2552
timestamp 1626908933
transform 1 0 14064 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2556
timestamp 1626908933
transform 1 0 14160 0 1 7659
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_248
timestamp 1626908933
transform 1 0 14400 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_849
timestamp 1626908933
transform 1 0 14400 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_697
timestamp 1626908933
transform 1 0 14352 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2664
timestamp 1626908933
transform 1 0 14352 0 1 8177
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_335
timestamp 1626908933
transform 1 0 14592 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_933
timestamp 1626908933
transform 1 0 14592 0 1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2578
timestamp 1626908933
transform 1 0 14736 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2577
timestamp 1626908933
transform 1 0 14736 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_611
timestamp 1626908933
transform 1 0 14736 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_610
timestamp 1626908933
transform 1 0 14736 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2563
timestamp 1626908933
transform 1 0 15024 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2562
timestamp 1626908933
transform 1 0 15024 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_596
timestamp 1626908933
transform 1 0 15024 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_595
timestamp 1626908933
transform 1 0 15024 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_619
timestamp 1626908933
transform 1 0 14976 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_262
timestamp 1626908933
transform 1 0 14976 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_92
timestamp 1626908933
transform 1 0 15072 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_31
timestamp 1626908933
transform 1 0 15072 0 1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2910
timestamp 1626908933
transform 1 0 15120 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_975
timestamp 1626908933
transform 1 0 15120 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2895
timestamp 1626908933
transform 1 0 15216 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2888
timestamp 1626908933
transform 1 0 15120 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_928
timestamp 1626908933
transform 1 0 15216 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_921
timestamp 1626908933
transform 1 0 15120 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_140
timestamp 1626908933
transform 1 0 15408 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2107
timestamp 1626908933
transform 1 0 15408 0 1 7881
box -32 -32 32 32
use L1M1_PR  L1M1_PR_978
timestamp 1626908933
transform 1 0 15312 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2913
timestamp 1626908933
transform 1 0 15312 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_139
timestamp 1626908933
transform 1 0 15408 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2106
timestamp 1626908933
transform 1 0 15408 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_157
timestamp 1626908933
transform 1 0 15312 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2092
timestamp 1626908933
transform 1 0 15312 0 1 8251
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_475
timestamp 1626908933
transform 1 0 15360 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1466
timestamp 1626908933
transform 1 0 15360 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_413
timestamp 1626908933
transform 1 0 15456 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1135
timestamp 1626908933
transform 1 0 15456 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_155
timestamp 1626908933
transform 1 0 15696 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2090
timestamp 1626908933
transform 1 0 15696 0 1 7881
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_498
timestamp 1626908933
transform 1 0 16100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1146
timestamp 1626908933
transform 1 0 16100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_498
timestamp 1626908933
transform 1 0 16100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1146
timestamp 1626908933
transform 1 0 16100 0 1 7992
box -100 -49 100 49
use M1M2_PR  M1M2_PR_594
timestamp 1626908933
transform 1 0 16272 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2561
timestamp 1626908933
transform 1 0 16272 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_602
timestamp 1626908933
transform 1 0 16272 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2537
timestamp 1626908933
transform 1 0 16272 0 1 8251
box -29 -23 29 23
use sky130_fd_sc_hs__nand4_1  sky130_fd_sc_hs__nand4_1_0
timestamp 1626908933
transform -1 0 16800 0 1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__nand4_1  sky130_fd_sc_hs__nand4_1_3
timestamp 1626908933
transform -1 0 16800 0 1 7992
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2654
timestamp 1626908933
transform 1 0 16560 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2651
timestamp 1626908933
transform 1 0 16368 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2089
timestamp 1626908933
transform 1 0 16464 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_719
timestamp 1626908933
transform 1 0 16560 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_716
timestamp 1626908933
transform 1 0 16368 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_154
timestamp 1626908933
transform 1 0 16464 0 1 7733
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2667
timestamp 1626908933
transform 1 0 16464 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_700
timestamp 1626908933
transform 1 0 16464 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2554
timestamp 1626908933
transform 1 0 16656 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1986
timestamp 1626908933
transform 1 0 16656 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_619
timestamp 1626908933
transform 1 0 16656 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_51
timestamp 1626908933
transform 1 0 16656 0 1 7733
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2013
timestamp 1626908933
transform 1 0 16656 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_46
timestamp 1626908933
transform 1 0 16656 0 1 7733
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1105
timestamp 1626908933
transform 1 0 16800 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_383
timestamp 1626908933
transform 1 0 16800 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_417
timestamp 1626908933
transform 1 0 17568 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1018
timestamp 1626908933
transform 1 0 17568 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_745
timestamp 1626908933
transform 1 0 17760 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1736
timestamp 1626908933
transform 1 0 17760 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_601
timestamp 1626908933
transform 1 0 17616 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2568
timestamp 1626908933
transform 1 0 17616 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_474
timestamp 1626908933
transform 1 0 18240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1465
timestamp 1626908933
transform 1 0 18240 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_687
timestamp 1626908933
transform 1 0 18096 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2654
timestamp 1626908933
transform 1 0 18096 0 1 8177
box -32 -32 32 32
use L1M1_PR  L1M1_PR_604
timestamp 1626908933
transform 1 0 18096 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_609
timestamp 1626908933
transform 1 0 17904 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2539
timestamp 1626908933
transform 1 0 18096 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2544
timestamp 1626908933
transform 1 0 17904 0 1 8251
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_4
timestamp 1626908933
transform -1 0 18240 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_66
timestamp 1626908933
transform -1 0 18240 0 1 7992
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_474
timestamp 1626908933
transform 1 0 18500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1122
timestamp 1626908933
transform 1 0 18500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_474
timestamp 1626908933
transform 1 0 18500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1122
timestamp 1626908933
transform 1 0 18500 0 1 7992
box -100 -49 100 49
use M1M2_PR  M1M2_PR_598
timestamp 1626908933
transform 1 0 18960 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_599
timestamp 1626908933
transform 1 0 18288 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2565
timestamp 1626908933
transform 1 0 18960 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2566
timestamp 1626908933
transform 1 0 18288 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_607
timestamp 1626908933
transform 1 0 18288 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2542
timestamp 1626908933
transform 1 0 18288 0 1 8251
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_78
timestamp 1626908933
transform 1 0 19104 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_9
timestamp 1626908933
transform 1 0 19104 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_338
timestamp 1626908933
transform 1 0 18336 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1060
timestamp 1626908933
transform 1 0 18336 0 1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_114
timestamp 1626908933
transform 1 0 19536 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2081
timestamp 1626908933
transform 1 0 19536 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_126
timestamp 1626908933
transform 1 0 19440 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2061
timestamp 1626908933
transform 1 0 19440 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_261
timestamp 1626908933
transform 1 0 19968 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_618
timestamp 1626908933
transform 1 0 19968 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_746
timestamp 1626908933
transform 1 0 20064 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1737
timestamp 1626908933
transform 1 0 20064 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_108
timestamp 1626908933
transform 1 0 20112 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2075
timestamp 1626908933
transform 1 0 20112 0 1 7733
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_222
timestamp 1626908933
transform 1 0 19584 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_820
timestamp 1626908933
transform 1 0 19584 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__maj3_1  sky130_fd_sc_hs__maj3_1_1
timestamp 1626908933
transform -1 0 20928 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__maj3_1  sky130_fd_sc_hs__maj3_1_3
timestamp 1626908933
transform -1 0 20928 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_122
timestamp 1626908933
transform 1 0 20304 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_709
timestamp 1626908933
transform 1 0 20400 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_943
timestamp 1626908933
transform 1 0 20496 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2057
timestamp 1626908933
transform 1 0 20304 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2644
timestamp 1626908933
transform 1 0 20400 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2878
timestamp 1626908933
transform 1 0 20496 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2639
timestamp 1626908933
transform 1 0 20688 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_704
timestamp 1626908933
transform 1 0 20688 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2858
timestamp 1626908933
transform 1 0 20688 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_891
timestamp 1626908933
transform 1 0 20688 0 1 7733
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1098
timestamp 1626908933
transform 1 0 20900 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_450
timestamp 1626908933
transform 1 0 20900 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1098
timestamp 1626908933
transform 1 0 20900 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_450
timestamp 1626908933
transform 1 0 20900 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1464
timestamp 1626908933
transform 1 0 20928 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_473
timestamp 1626908933
transform 1 0 20928 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_286
timestamp 1626908933
transform 1 0 21024 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1008
timestamp 1626908933
transform 1 0 21024 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2477
timestamp 1626908933
transform 1 0 21456 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_542
timestamp 1626908933
transform 1 0 21456 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2479
timestamp 1626908933
transform 1 0 21648 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2474
timestamp 1626908933
transform 1 0 21744 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_544
timestamp 1626908933
transform 1 0 21648 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_539
timestamp 1626908933
transform 1 0 21744 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2509
timestamp 1626908933
transform 1 0 21648 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_542
timestamp 1626908933
transform 1 0 21648 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2503
timestamp 1626908933
transform 1 0 21840 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_536
timestamp 1626908933
transform 1 0 21840 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2500
timestamp 1626908933
transform 1 0 21072 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_533
timestamp 1626908933
transform 1 0 21072 0 1 7807
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2469
timestamp 1626908933
transform 1 0 21552 0 1 7807
box -29 -23 29 23
use L1M1_PR  L1M1_PR_534
timestamp 1626908933
transform 1 0 21552 0 1 7807
box -29 -23 29 23
use M1M2_PR  M1M2_PR_95
timestamp 1626908933
transform 1 0 21456 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2062
timestamp 1626908933
transform 1 0 21456 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_550
timestamp 1626908933
transform 1 0 21744 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2485
timestamp 1626908933
transform 1 0 21744 0 1 8177
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_11
timestamp 1626908933
transform 1 0 21792 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_73
timestamp 1626908933
transform 1 0 21792 0 1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2472
timestamp 1626908933
transform 1 0 21936 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2042
timestamp 1626908933
transform 1 0 21936 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_537
timestamp 1626908933
transform 1 0 21936 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_107
timestamp 1626908933
transform 1 0 21936 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2476
timestamp 1626908933
transform 1 0 22224 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_541
timestamp 1626908933
transform 1 0 22224 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2507
timestamp 1626908933
transform 1 0 22128 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2506
timestamp 1626908933
transform 1 0 22128 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_540
timestamp 1626908933
transform 1 0 22128 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_539
timestamp 1626908933
transform 1 0 22128 0 1 8103
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1463
timestamp 1626908933
transform 1 0 22368 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_472
timestamp 1626908933
transform 1 0 22368 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_848
timestamp 1626908933
transform 1 0 22176 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_247
timestamp 1626908933
transform 1 0 22176 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_534
timestamp 1626908933
transform 1 0 22800 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2501
timestamp 1626908933
transform 1 0 22800 0 1 7659
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_255
timestamp 1626908933
transform 1 0 22464 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_977
timestamp 1626908933
transform 1 0 22464 0 1 7992
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_426
timestamp 1626908933
transform 1 0 23300 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1074
timestamp 1626908933
transform 1 0 23300 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_426
timestamp 1626908933
transform 1 0 23300 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1074
timestamp 1626908933
transform 1 0 23300 0 1 7992
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2543
timestamp 1626908933
transform 1 0 22992 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_576
timestamp 1626908933
transform 1 0 22992 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2517
timestamp 1626908933
transform 1 0 23280 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_582
timestamp 1626908933
transform 1 0 23280 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2511
timestamp 1626908933
transform 1 0 23376 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_576
timestamp 1626908933
transform 1 0 23376 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2679
timestamp 1626908933
transform 1 0 23568 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_744
timestamp 1626908933
transform 1 0 23568 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2687
timestamp 1626908933
transform 1 0 23568 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_720
timestamp 1626908933
transform 1 0 23568 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_161
timestamp 1626908933
transform 1 0 23616 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_759
timestamp 1626908933
transform 1 0 23616 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_2
timestamp 1626908933
transform -1 0 23616 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_10
timestamp 1626908933
transform -1 0 23616 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_418
timestamp 1626908933
transform 1 0 24000 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1019
timestamp 1626908933
transform 1 0 24000 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_747
timestamp 1626908933
transform 1 0 24192 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1738
timestamp 1626908933
transform 1 0 24192 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_13
timestamp 1626908933
transform -1 0 24576 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_74
timestamp 1626908933
transform -1 0 24576 0 1 7992
box -38 -49 326 715
use M1M2_PR  M1M2_PR_882
timestamp 1626908933
transform 1 0 24240 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2849
timestamp 1626908933
transform 1 0 24240 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_930
timestamp 1626908933
transform 1 0 24336 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2865
timestamp 1626908933
transform 1 0 24336 0 1 8103
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_20
timestamp 1626908933
transform 1 0 24576 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_72
timestamp 1626908933
transform 1 0 24576 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_260
timestamp 1626908933
transform 1 0 24960 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_617
timestamp 1626908933
transform 1 0 24960 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_419
timestamp 1626908933
transform 1 0 25056 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1020
timestamp 1626908933
transform 1 0 25056 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_748
timestamp 1626908933
transform 1 0 25248 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1739
timestamp 1626908933
transform 1 0 25248 0 1 7992
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1050
timestamp 1626908933
transform 1 0 25700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_402
timestamp 1626908933
transform 1 0 25700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1050
timestamp 1626908933
transform 1 0 25700 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_402
timestamp 1626908933
transform 1 0 25700 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3515
timestamp 1626908933
transform 1 0 25392 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1580
timestamp 1626908933
transform 1 0 25392 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3459
timestamp 1626908933
transform 1 0 25488 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1492
timestamp 1626908933
transform 1 0 25488 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2933
timestamp 1626908933
transform 1 0 25488 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_966
timestamp 1626908933
transform 1 0 25488 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2963
timestamp 1626908933
transform 1 0 25584 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1028
timestamp 1626908933
transform 1 0 25584 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_21
timestamp 1626908933
transform 1 0 25344 0 1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_60
timestamp 1626908933
transform 1 0 25344 0 1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_847
timestamp 1626908933
transform 1 0 25920 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_246
timestamp 1626908933
transform 1 0 25920 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_706
timestamp 1626908933
transform 1 0 26112 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_108
timestamp 1626908933
transform 1 0 26112 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_885
timestamp 1626908933
transform 1 0 26496 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_163
timestamp 1626908933
transform 1 0 26496 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_686
timestamp 1626908933
transform 1 0 27264 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_88
timestamp 1626908933
transform 1 0 27264 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_852
timestamp 1626908933
transform 1 0 27648 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_130
timestamp 1626908933
transform 1 0 27648 0 1 7992
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1026
timestamp 1626908933
transform 1 0 28100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_378
timestamp 1626908933
transform 1 0 28100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1026
timestamp 1626908933
transform 1 0 28100 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_378
timestamp 1626908933
transform 1 0 28100 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_11
timestamp 1626908933
transform 1 0 28416 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_80
timestamp 1626908933
transform 1 0 28416 0 1 7992
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2482
timestamp 1626908933
transform 1 0 28560 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_547
timestamp 1626908933
transform 1 0 28560 0 1 8177
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1462
timestamp 1626908933
transform 1 0 28896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_471
timestamp 1626908933
transform 1 0 28896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_817
timestamp 1626908933
transform 1 0 28992 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_95
timestamp 1626908933
transform 1 0 28992 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1740
timestamp 1626908933
transform 1 0 29856 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1461
timestamp 1626908933
transform 1 0 29760 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_749
timestamp 1626908933
transform 1 0 29856 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_470
timestamp 1626908933
transform 1 0 29760 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_846
timestamp 1626908933
transform 1 0 30048 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_245
timestamp 1626908933
transform 1 0 30048 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_616
timestamp 1626908933
transform 1 0 29952 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_259
timestamp 1626908933
transform 1 0 29952 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1460
timestamp 1626908933
transform 1 0 30240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_469
timestamp 1626908933
transform 1 0 30240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_778
timestamp 1626908933
transform 1 0 30336 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_56
timestamp 1626908933
transform 1 0 30336 0 1 7992
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1002
timestamp 1626908933
transform 1 0 30500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_354
timestamp 1626908933
transform 1 0 30500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1002
timestamp 1626908933
transform 1 0 30500 0 1 7992
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_354
timestamp 1626908933
transform 1 0 30500 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1459
timestamp 1626908933
transform 1 0 31104 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_468
timestamp 1626908933
transform 1 0 31104 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_739
timestamp 1626908933
transform 1 0 31200 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_17
timestamp 1626908933
transform 1 0 31200 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1741
timestamp 1626908933
transform 1 0 31968 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_750
timestamp 1626908933
transform 1 0 31968 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3887
timestamp 1626908933
transform 1 0 144 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1920
timestamp 1626908933
transform 1 0 144 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1458
timestamp 1626908933
transform 1 0 0 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_467
timestamp 1626908933
transform 1 0 0 0 -1 9324
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_977
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_329
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_977
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_329
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1195
timestamp 1626908933
transform 1 0 96 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_597
timestamp 1626908933
transform 1 0 96 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_466
timestamp 1626908933
transform 1 0 480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_751
timestamp 1626908933
transform 1 0 576 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1457
timestamp 1626908933
transform 1 0 480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1742
timestamp 1626908933
transform 1 0 576 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1287
timestamp 1626908933
transform 1 0 912 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1889
timestamp 1626908933
transform 1 0 720 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3222
timestamp 1626908933
transform 1 0 912 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3824
timestamp 1626908933
transform 1 0 720 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_1
timestamp 1626908933
transform 1 0 672 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_6
timestamp 1626908933
transform 1 0 672 0 -1 9324
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1138
timestamp 1626908933
transform 1 0 1392 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1756
timestamp 1626908933
transform 1 0 1200 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3105
timestamp 1626908933
transform 1 0 1392 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3723
timestamp 1626908933
transform 1 0 1200 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_335
timestamp 1626908933
transform 1 0 1776 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2270
timestamp 1626908933
transform 1 0 1776 0 1 8399
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1215
timestamp 1626908933
transform 1 0 1488 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1919
timestamp 1626908933
transform 1 0 1008 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3182
timestamp 1626908933
transform 1 0 1488 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3886
timestamp 1626908933
transform 1 0 1008 0 1 9065
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_683
timestamp 1626908933
transform 1 0 1152 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1405
timestamp 1626908933
transform 1 0 1152 0 -1 9324
box -38 -49 806 715
use M1M2_PR  M1M2_PR_311
timestamp 1626908933
transform 1 0 2256 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2278
timestamp 1626908933
transform 1 0 2256 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1887
timestamp 1626908933
transform 1 0 1968 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3822
timestamp 1626908933
transform 1 0 1968 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3342
timestamp 1626908933
transform 1 0 2352 0 1 8473
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1407
timestamp 1626908933
transform 1 0 2352 0 1 8473
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1743
timestamp 1626908933
transform 1 0 2400 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_752
timestamp 1626908933
transform 1 0 2400 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_615
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_258
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3821
timestamp 1626908933
transform 1 0 2640 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3701
timestamp 1626908933
transform 1 0 2544 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1886
timestamp 1626908933
transform 1 0 2640 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1766
timestamp 1626908933
transform 1 0 2544 0 1 8547
box -29 -23 29 23
use sky130_fd_sc_hs__nand3b_2  sky130_fd_sc_hs__nand3b_2_0
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand3b_2  sky130_fd_sc_hs__nand3b_2_1
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nor2_2  sky130_fd_sc_hs__nor2_2_1
timestamp 1626908933
transform 1 0 1920 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nor2_2  sky130_fd_sc_hs__nor2_2_3
timestamp 1626908933
transform 1 0 1920 0 -1 9324
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1205
timestamp 1626908933
transform 1 0 3600 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3140
timestamp 1626908933
transform 1 0 3600 0 1 8769
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_305
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_953
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_305
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_953
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3721
timestamp 1626908933
transform 1 0 2928 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1786
timestamp 1626908933
transform 1 0 2928 0 1 8917
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3738
timestamp 1626908933
transform 1 0 2928 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1771
timestamp 1626908933
transform 1 0 2928 0 1 8917
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3631
timestamp 1626908933
transform 1 0 2832 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1696
timestamp 1626908933
transform 1 0 2832 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3719
timestamp 1626908933
transform 1 0 3120 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1752
timestamp 1626908933
transform 1 0 3120 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3697
timestamp 1626908933
transform 1 0 3216 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1762
timestamp 1626908933
transform 1 0 3216 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3567
timestamp 1626908933
transform 1 0 3504 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1600
timestamp 1626908933
transform 1 0 3504 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3628
timestamp 1626908933
transform 1 0 3600 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1693
timestamp 1626908933
transform 1 0 3600 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_129
timestamp 1626908933
transform -1 0 3936 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_60
timestamp 1626908933
transform -1 0 3936 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_753
timestamp 1626908933
transform 1 0 3936 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1744
timestamp 1626908933
transform 1 0 3936 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1153
timestamp 1626908933
transform 1 0 3792 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3120
timestamp 1626908933
transform 1 0 3792 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1882
timestamp 1626908933
transform 1 0 3984 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1883
timestamp 1626908933
transform 1 0 3984 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3817
timestamp 1626908933
transform 1 0 3984 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3818
timestamp 1626908933
transform 1 0 3984 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1139
timestamp 1626908933
transform 1 0 4176 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1326
timestamp 1626908933
transform 1 0 4368 0 1 8473
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3106
timestamp 1626908933
transform 1 0 4176 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3293
timestamp 1626908933
transform 1 0 4368 0 1 8473
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1209
timestamp 1626908933
transform 1 0 4176 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1775
timestamp 1626908933
transform 1 0 4272 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3144
timestamp 1626908933
transform 1 0 4176 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3710
timestamp 1626908933
transform 1 0 4272 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_3
timestamp 1626908933
transform 1 0 4032 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_8
timestamp 1626908933
transform 1 0 4032 0 -1 9324
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3157
timestamp 1626908933
transform 1 0 4656 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1222
timestamp 1626908933
transform 1 0 4656 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3709
timestamp 1626908933
transform 1 0 4656 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1774
timestamp 1626908933
transform 1 0 4656 0 1 8917
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3102
timestamp 1626908933
transform 1 0 4848 0 1 8843
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1135
timestamp 1626908933
transform 1 0 4848 0 1 8843
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3147
timestamp 1626908933
transform 1 0 4560 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1212
timestamp 1626908933
transform 1 0 4560 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3109
timestamp 1626908933
transform 1 0 4560 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1142
timestamp 1626908933
transform 1 0 4560 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3814
timestamp 1626908933
transform 1 0 4752 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1879
timestamp 1626908933
transform 1 0 4752 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3101
timestamp 1626908933
transform 1 0 4848 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1134
timestamp 1626908933
transform 1 0 4848 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3139
timestamp 1626908933
transform 1 0 4848 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1204
timestamp 1626908933
transform 1 0 4848 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3712
timestamp 1626908933
transform 1 0 4464 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1777
timestamp 1626908933
transform 1 0 4464 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3711
timestamp 1626908933
transform 1 0 4944 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1776
timestamp 1626908933
transform 1 0 4944 0 1 8991
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_929
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_281
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_929
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_281
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3345
timestamp 1626908933
transform 1 0 5232 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1410
timestamp 1626908933
transform 1 0 5232 0 1 9139
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1456
timestamp 1626908933
transform 1 0 5184 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_465
timestamp 1626908933
transform 1 0 5184 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_120
timestamp 1626908933
transform 1 0 4896 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_58
timestamp 1626908933
transform 1 0 4896 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_606
timestamp 1626908933
transform 1 0 5280 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1328
timestamp 1626908933
transform 1 0 5280 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_7
timestamp 1626908933
transform 1 0 4512 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_15
timestamp 1626908933
transform 1 0 4512 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nor2b_2  sky130_fd_sc_hs__nor2b_2_1
timestamp 1626908933
transform -1 0 6720 0 -1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__nor2b_2  sky130_fd_sc_hs__nor2b_2_0
timestamp 1626908933
transform -1 0 6720 0 -1 9324
box -38 -49 710 715
use L1M1_PR  L1M1_PR_3811
timestamp 1626908933
transform 1 0 6192 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1876
timestamp 1626908933
transform 1 0 6192 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1328
timestamp 1626908933
transform 1 0 6480 0 1 9139
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3295
timestamp 1626908933
transform 1 0 6480 0 1 9139
box -32 -32 32 32
use L1M1_PR  L1M1_PR_398
timestamp 1626908933
transform 1 0 6576 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2333
timestamp 1626908933
transform 1 0 6576 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2332
timestamp 1626908933
transform 1 0 6768 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_397
timestamp 1626908933
transform 1 0 6768 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2342
timestamp 1626908933
transform 1 0 6672 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_375
timestamp 1626908933
transform 1 0 6672 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2068
timestamp 1626908933
transform 1 0 6960 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_133
timestamp 1626908933
transform 1 0 6960 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2341
timestamp 1626908933
transform 1 0 6672 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2089
timestamp 1626908933
transform 1 0 6864 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_374
timestamp 1626908933
transform 1 0 6672 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_122
timestamp 1626908933
transform 1 0 6864 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1021
timestamp 1626908933
transform 1 0 6720 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_420
timestamp 1626908933
transform 1 0 6720 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_12
timestamp 1626908933
transform -1 0 7488 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_51
timestamp 1626908933
transform -1 0 7488 0 -1 9324
box -38 -49 614 715
use M1M2_PR  M1M2_PR_904
timestamp 1626908933
transform 1 0 7056 0 1 9139
box -32 -32 32 32
use M1M2_PR  M1M2_PR_907
timestamp 1626908933
transform 1 0 7248 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2871
timestamp 1626908933
transform 1 0 7056 0 1 9139
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2874
timestamp 1626908933
transform 1 0 7248 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_953
timestamp 1626908933
transform 1 0 7056 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_956
timestamp 1626908933
transform 1 0 7248 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2888
timestamp 1626908933
transform 1 0 7056 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2891
timestamp 1626908933
transform 1 0 7248 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_257
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_614
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_257
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_905
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_257
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_905
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_471
timestamp 1626908933
transform 1 0 7584 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1069
timestamp 1626908933
transform 1 0 7584 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_39
timestamp 1626908933
transform 1 0 8064 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_0
timestamp 1626908933
transform 1 0 8064 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1745
timestamp 1626908933
transform 1 0 7968 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_754
timestamp 1626908933
transform 1 0 7968 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_25
timestamp 1626908933
transform 1 0 8592 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_843
timestamp 1626908933
transform 1 0 8496 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_847
timestamp 1626908933
transform 1 0 8304 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1960
timestamp 1626908933
transform 1 0 8592 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2778
timestamp 1626908933
transform 1 0 8496 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2782
timestamp 1626908933
transform 1 0 8304 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_464
timestamp 1626908933
transform 1 0 8640 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1455
timestamp 1626908933
transform 1 0 8640 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_447
timestamp 1626908933
transform 1 0 8736 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1045
timestamp 1626908933
transform 1 0 8736 0 -1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2779
timestamp 1626908933
transform 1 0 8976 0 1 8843
box -32 -32 32 32
use M1M2_PR  M1M2_PR_812
timestamp 1626908933
transform 1 0 8976 0 1 8843
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2780
timestamp 1626908933
transform 1 0 9264 0 1 8843
box -29 -23 29 23
use L1M1_PR  L1M1_PR_845
timestamp 1626908933
transform 1 0 9264 0 1 8843
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1989
timestamp 1626908933
transform 1 0 9072 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_22
timestamp 1626908933
transform 1 0 9072 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2774
timestamp 1626908933
transform 1 0 9168 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_807
timestamp 1626908933
transform 1 0 9168 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2776
timestamp 1626908933
transform 1 0 9168 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_841
timestamp 1626908933
transform 1 0 9168 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1958
timestamp 1626908933
transform 1 0 9360 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_23
timestamp 1626908933
transform 1 0 9360 0 1 9065
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_22
timestamp 1626908933
transform 1 0 9120 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_83
timestamp 1626908933
transform 1 0 9120 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_436
timestamp 1626908933
transform 1 0 9408 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1034
timestamp 1626908933
transform 1 0 9408 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_421
timestamp 1626908933
transform 1 0 9792 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1022
timestamp 1626908933
transform 1 0 9792 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_704
timestamp 1626908933
transform 1 0 9648 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2671
timestamp 1626908933
transform 1 0 9648 0 1 8917
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_755
timestamp 1626908933
transform 1 0 9984 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1746
timestamp 1626908933
transform 1 0 9984 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_21
timestamp 1626908933
transform 1 0 10128 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1956
timestamp 1626908933
transform 1 0 10128 0 1 8991
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_233
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_881
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_233
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_881
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_2
timestamp 1626908933
transform -1 0 10656 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_8
timestamp 1626908933
transform -1 0 10656 0 -1 9324
box -38 -49 614 715
use M1M2_PR  M1M2_PR_2734
timestamp 1626908933
transform 1 0 10320 0 1 8473
box -32 -32 32 32
use M1M2_PR  M1M2_PR_767
timestamp 1626908933
transform 1 0 10320 0 1 8473
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2731
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2659
timestamp 1626908933
transform 1 0 10416 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_796
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_724
timestamp 1626908933
transform 1 0 10416 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2733
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_766
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2585
timestamp 1626908933
transform 1 0 10512 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_650
timestamp 1626908933
transform 1 0 10512 0 1 9139
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_244
timestamp 1626908933
transform 1 0 10656 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_845
timestamp 1626908933
transform 1 0 10656 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_18
timestamp 1626908933
transform 1 0 10608 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1985
timestamp 1626908933
transform 1 0 10608 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_17
timestamp 1626908933
transform 1 0 10608 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1952
timestamp 1626908933
transform 1 0 10608 0 1 9065
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_463
timestamp 1626908933
transform 1 0 10848 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1454
timestamp 1626908933
transform 1 0 10848 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2602
timestamp 1626908933
transform 1 0 10992 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_635
timestamp 1626908933
transform 1 0 10992 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1004
timestamp 1626908933
transform 1 0 10944 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_406
timestamp 1626908933
transform 1 0 10944 0 -1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_643
timestamp 1626908933
transform 1 0 11376 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2578
timestamp 1626908933
transform 1 0 11376 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_632
timestamp 1626908933
transform 1 0 11568 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2599
timestamp 1626908933
transform 1 0 11568 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_640
timestamp 1626908933
transform 1 0 11568 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2575
timestamp 1626908933
transform 1 0 11568 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_637
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2604
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_646
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2581
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_633
timestamp 1626908933
transform 1 0 11760 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2568
timestamp 1626908933
transform 1 0 11760 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_649
timestamp 1626908933
transform 1 0 11856 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2584
timestamp 1626908933
transform 1 0 11856 0 1 9065
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_844
timestamp 1626908933
transform 1 0 11904 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_243
timestamp 1626908933
transform 1 0 11904 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_2
timestamp 1626908933
transform -1 0 11904 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_15
timestamp 1626908933
transform -1 0 11904 0 -1 9324
box -38 -49 614 715
use M1M2_PR  M1M2_PR_622
timestamp 1626908933
transform 1 0 11952 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_639
timestamp 1626908933
transform 1 0 12144 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_640
timestamp 1626908933
transform 1 0 12144 0 1 8473
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2589
timestamp 1626908933
transform 1 0 11952 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2606
timestamp 1626908933
transform 1 0 12144 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2607
timestamp 1626908933
transform 1 0 12144 0 1 8473
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_256
timestamp 1626908933
transform 1 0 12480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_613
timestamp 1626908933
transform 1 0 12480 0 -1 9324
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_209
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_857
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_209
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_857
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_365
timestamp 1626908933
transform 1 0 12576 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_381
timestamp 1626908933
transform 1 0 12096 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_963
timestamp 1626908933
transform 1 0 12576 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_979
timestamp 1626908933
transform 1 0 12096 0 -1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2726
timestamp 1626908933
transform 1 0 12816 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_791
timestamp 1626908933
transform 1 0 12816 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2728
timestamp 1626908933
transform 1 0 12816 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_761
timestamp 1626908933
transform 1 0 12816 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2622
timestamp 1626908933
transform 1 0 13200 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2583
timestamp 1626908933
transform 1 0 13104 0 1 8473
box -29 -23 29 23
use L1M1_PR  L1M1_PR_687
timestamp 1626908933
transform 1 0 13200 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_648
timestamp 1626908933
transform 1 0 13104 0 1 8473
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2637
timestamp 1626908933
transform 1 0 13200 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_670
timestamp 1626908933
transform 1 0 13200 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_463
timestamp 1626908933
transform 1 0 12960 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1185
timestamp 1626908933
transform 1 0 12960 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1023
timestamp 1626908933
transform 1 0 13728 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_422
timestamp 1626908933
transform 1 0 13728 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_756
timestamp 1626908933
transform 1 0 13920 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1747
timestamp 1626908933
transform 1 0 13920 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_982
timestamp 1626908933
transform 1 0 13968 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2917
timestamp 1626908933
transform 1 0 13968 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_769
timestamp 1626908933
transform 1 0 14256 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2704
timestamp 1626908933
transform 1 0 14256 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_7
timestamp 1626908933
transform 1 0 14400 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_30
timestamp 1626908933
transform 1 0 14400 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_29
timestamp 1626908933
transform -1 0 14400 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_91
timestamp 1626908933
transform -1 0 14400 0 -1 9324
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_185
timestamp 1626908933
transform 1 0 14900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_833
timestamp 1626908933
transform 1 0 14900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_185
timestamp 1626908933
transform 1 0 14900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_833
timestamp 1626908933
transform 1 0 14900 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1748
timestamp 1626908933
transform 1 0 15168 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_757
timestamp 1626908933
transform 1 0 15168 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_927
timestamp 1626908933
transform 1 0 15216 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2894
timestamp 1626908933
transform 1 0 15216 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_980
timestamp 1626908933
transform 1 0 15216 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2915
timestamp 1626908933
transform 1 0 15216 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_981
timestamp 1626908933
transform 1 0 15312 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2916
timestamp 1626908933
transform 1 0 15312 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_926
timestamp 1626908933
transform 1 0 15216 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2893
timestamp 1626908933
transform 1 0 15216 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_979
timestamp 1626908933
transform 1 0 15216 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2914
timestamp 1626908933
transform 1 0 15216 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_744
timestamp 1626908933
transform 1 0 15312 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2711
timestamp 1626908933
transform 1 0 15312 0 1 9065
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_97
timestamp 1626908933
transform -1 0 15552 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_35
timestamp 1626908933
transform -1 0 15552 0 -1 9324
box -38 -49 326 715
use L1M1_PR  L1M1_PR_767
timestamp 1626908933
transform 1 0 15504 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2702
timestamp 1626908933
transform 1 0 15504 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1982
timestamp 1626908933
transform 1 0 15600 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_15
timestamp 1626908933
transform 1 0 15600 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1749
timestamp 1626908933
transform 1 0 16320 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_758
timestamp 1626908933
transform 1 0 16320 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1134
timestamp 1626908933
transform 1 0 15552 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_412
timestamp 1626908933
transform 1 0 15552 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__a211oi_1  sky130_fd_sc_hs__a211oi_1_2
timestamp 1626908933
transform 1 0 16416 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__a211oi_1  sky130_fd_sc_hs__a211oi_1_0
timestamp 1626908933
transform 1 0 16416 0 -1 9324
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2658
timestamp 1626908933
transform 1 0 16368 0 1 8843
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2650
timestamp 1626908933
transform 1 0 16368 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_723
timestamp 1626908933
transform 1 0 16368 0 1 8843
box -29 -23 29 23
use L1M1_PR  L1M1_PR_715
timestamp 1626908933
transform 1 0 16368 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2666
timestamp 1626908933
transform 1 0 16464 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_699
timestamp 1626908933
transform 1 0 16464 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_696
timestamp 1626908933
transform 1 0 16848 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2663
timestamp 1626908933
transform 1 0 16848 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_16
timestamp 1626908933
transform 1 0 16656 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_718
timestamp 1626908933
transform 1 0 16848 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_729
timestamp 1626908933
transform 1 0 16752 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1951
timestamp 1626908933
transform 1 0 16656 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2653
timestamp 1626908933
transform 1 0 16848 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2664
timestamp 1626908933
transform 1 0 16752 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_462
timestamp 1626908933
transform 1 0 16992 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1453
timestamp 1626908933
transform 1 0 16992 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_731
timestamp 1626908933
transform 1 0 16944 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2666
timestamp 1626908933
transform 1 0 16944 0 1 9065
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_161
timestamp 1626908933
transform 1 0 17300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_809
timestamp 1626908933
transform 1 0 17300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_161
timestamp 1626908933
transform 1 0 17300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_809
timestamp 1626908933
transform 1 0 17300 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_282
timestamp 1626908933
transform 1 0 17088 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_880
timestamp 1626908933
transform 1 0 17088 0 -1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2676
timestamp 1626908933
transform 1 0 17328 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2556
timestamp 1626908933
transform 1 0 17520 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_709
timestamp 1626908933
transform 1 0 17328 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_589
timestamp 1626908933
transform 1 0 17520 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_869
timestamp 1626908933
transform 1 0 17568 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_271
timestamp 1626908933
transform 1 0 17568 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_612
timestamp 1626908933
transform 1 0 17472 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_255
timestamp 1626908933
transform 1 0 17472 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2531
timestamp 1626908933
transform 1 0 17904 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_596
timestamp 1626908933
transform 1 0 17904 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2653
timestamp 1626908933
transform 1 0 18096 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_686
timestamp 1626908933
transform 1 0 18096 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2752
timestamp 1626908933
transform 1 0 18000 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_785
timestamp 1626908933
transform 1 0 18000 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2750
timestamp 1626908933
transform 1 0 18096 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2580
timestamp 1626908933
transform 1 0 18192 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_815
timestamp 1626908933
transform 1 0 18096 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_645
timestamp 1626908933
transform 1 0 18192 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2640
timestamp 1626908933
transform 1 0 18384 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_705
timestamp 1626908933
transform 1 0 18384 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2080
timestamp 1626908933
transform 1 0 18480 0 1 8473
box -32 -32 32 32
use M1M2_PR  M1M2_PR_113
timestamp 1626908933
transform 1 0 18480 0 1 8473
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2060
timestamp 1626908933
transform 1 0 18480 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_125
timestamp 1626908933
transform 1 0 18480 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2079
timestamp 1626908933
transform 1 0 18480 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_112
timestamp 1626908933
transform 1 0 18480 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_843
timestamp 1626908933
transform 1 0 18528 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_242
timestamp 1626908933
transform 1 0 18528 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_2
timestamp 1626908933
transform -1 0 18528 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_8
timestamp 1626908933
transform -1 0 18528 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1452
timestamp 1626908933
transform 1 0 18720 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_461
timestamp 1626908933
transform 1 0 18720 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_844
timestamp 1626908933
transform 1 0 18816 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_246
timestamp 1626908933
transform 1 0 18816 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_68
timestamp 1626908933
transform -1 0 19488 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_7
timestamp 1626908933
transform -1 0 19488 0 -1 9324
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2147
timestamp 1626908933
transform 1 0 19248 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_212
timestamp 1626908933
transform 1 0 19248 0 1 9065
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2159
timestamp 1626908933
transform 1 0 19248 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_192
timestamp 1626908933
transform 1 0 19248 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2058
timestamp 1626908933
transform 1 0 20112 0 1 8473
box -29 -23 29 23
use L1M1_PR  L1M1_PR_123
timestamp 1626908933
transform 1 0 20112 0 1 8473
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2074
timestamp 1626908933
transform 1 0 20112 0 1 8473
box -32 -32 32 32
use M1M2_PR  M1M2_PR_107
timestamp 1626908933
transform 1 0 20112 0 1 8473
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2693
timestamp 1626908933
transform 1 0 19440 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_758
timestamp 1626908933
transform 1 0 19440 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2702
timestamp 1626908933
transform 1 0 19536 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_735
timestamp 1626908933
transform 1 0 19536 0 1 8547
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_785
timestamp 1626908933
transform 1 0 19700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_137
timestamp 1626908933
transform 1 0 19700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_785
timestamp 1626908933
transform 1 0 19700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_137
timestamp 1626908933
transform 1 0 19700 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2692
timestamp 1626908933
transform 1 0 19536 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_757
timestamp 1626908933
transform 1 0 19536 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2701
timestamp 1626908933
transform 1 0 19536 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_734
timestamp 1626908933
transform 1 0 19536 0 1 8769
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_8
timestamp 1626908933
transform 1 0 19488 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_31
timestamp 1626908933
transform 1 0 19488 0 -1 9324
box -38 -49 806 715
use M1M2_PR  M1M2_PR_523
timestamp 1626908933
transform 1 0 20688 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_691
timestamp 1626908933
transform 1 0 20496 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2490
timestamp 1626908933
transform 1 0 20688 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2658
timestamp 1626908933
transform 1 0 20496 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_520
timestamp 1626908933
transform 1 0 20880 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2455
timestamp 1626908933
transform 1 0 20880 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2663
timestamp 1626908933
transform 1 0 20304 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_728
timestamp 1626908933
transform 1 0 20304 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2459
timestamp 1626908933
transform 1 0 20400 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_524
timestamp 1626908933
transform 1 0 20400 0 1 9065
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2657
timestamp 1626908933
transform 1 0 20496 0 1 9139
box -32 -32 32 32
use M1M2_PR  M1M2_PR_690
timestamp 1626908933
transform 1 0 20496 0 1 9139
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2486
timestamp 1626908933
transform 1 0 20688 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_551
timestamp 1626908933
transform 1 0 20688 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2643
timestamp 1626908933
transform 1 0 20496 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_708
timestamp 1626908933
transform 1 0 20496 0 1 9139
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_9
timestamp 1626908933
transform 1 0 20832 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_32
timestamp 1626908933
transform 1 0 20832 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_1
timestamp 1626908933
transform -1 0 20832 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_7
timestamp 1626908933
transform -1 0 20832 0 -1 9324
box -38 -49 614 715
use M1M2_PR  M1M2_PR_541
timestamp 1626908933
transform 1 0 21648 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_546
timestamp 1626908933
transform 1 0 21744 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2508
timestamp 1626908933
transform 1 0 21648 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2513
timestamp 1626908933
transform 1 0 21744 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_543
timestamp 1626908933
transform 1 0 21648 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_549
timestamp 1626908933
transform 1 0 21744 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2478
timestamp 1626908933
transform 1 0 21648 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2484
timestamp 1626908933
transform 1 0 21744 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_545
timestamp 1626908933
transform 1 0 21744 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2512
timestamp 1626908933
transform 1 0 21744 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_546
timestamp 1626908933
transform 1 0 21840 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2481
timestamp 1626908933
transform 1 0 21840 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__maj3_1  sky130_fd_sc_hs__maj3_1_0
timestamp 1626908933
transform 1 0 21600 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__maj3_1  sky130_fd_sc_hs__maj3_1_2
timestamp 1626908933
transform 1 0 21600 0 -1 9324
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_761
timestamp 1626908933
transform 1 0 22100 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_113
timestamp 1626908933
transform 1 0 22100 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_761
timestamp 1626908933
transform 1 0 22100 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_113
timestamp 1626908933
transform 1 0 22100 0 1 8658
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2757
timestamp 1626908933
transform 1 0 21936 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_790
timestamp 1626908933
transform 1 0 21936 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2757
timestamp 1626908933
transform 1 0 22128 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2483
timestamp 1626908933
transform 1 0 22128 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_822
timestamp 1626908933
transform 1 0 22128 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_548
timestamp 1626908933
transform 1 0 22128 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2679
timestamp 1626908933
transform 1 0 22320 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_712
timestamp 1626908933
transform 1 0 22320 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1750
timestamp 1626908933
transform 1 0 22368 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_759
timestamp 1626908933
transform 1 0 22368 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_611
timestamp 1626908933
transform 1 0 22464 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_254
timestamp 1626908933
transform 1 0 22464 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_254
timestamp 1626908933
transform 1 0 22560 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_976
timestamp 1626908933
transform 1 0 22560 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_760
timestamp 1626908933
transform 1 0 23328 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1751
timestamp 1626908933
transform 1 0 23328 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_544
timestamp 1626908933
transform 1 0 23088 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2511
timestamp 1626908933
transform 1 0 23088 0 1 8917
box -32 -32 32 32
use L1M1_PR  L1M1_PR_734
timestamp 1626908933
transform 1 0 23280 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2669
timestamp 1626908933
transform 1 0 23280 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2678
timestamp 1626908933
transform 1 0 23568 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_743
timestamp 1626908933
transform 1 0 23568 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2686
timestamp 1626908933
transform 1 0 23568 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2538
timestamp 1626908933
transform 1 0 23472 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_719
timestamp 1626908933
transform 1 0 23568 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_571
timestamp 1626908933
transform 1 0 23472 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2500
timestamp 1626908933
transform 1 0 23664 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2029
timestamp 1626908933
transform 1 0 23472 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_565
timestamp 1626908933
transform 1 0 23664 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_94
timestamp 1626908933
transform 1 0 23472 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2527
timestamp 1626908933
transform 1 0 23664 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_560
timestamp 1626908933
transform 1 0 23664 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_67
timestamp 1626908933
transform 1 0 23424 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_5
timestamp 1626908933
transform 1 0 23424 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_241
timestamp 1626908933
transform 1 0 23712 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_842
timestamp 1626908933
transform 1 0 23712 0 -1 9324
box -38 -49 230 715
use L1M1_PR  L1M1_PR_105
timestamp 1626908933
transform 1 0 24240 0 1 8473
box -29 -23 29 23
use L1M1_PR  L1M1_PR_928
timestamp 1626908933
transform 1 0 24624 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2040
timestamp 1626908933
transform 1 0 24240 0 1 8473
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2863
timestamp 1626908933
transform 1 0 24624 0 1 8547
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_89
timestamp 1626908933
transform 1 0 24500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_737
timestamp 1626908933
transform 1 0 24500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_89
timestamp 1626908933
transform 1 0 24500 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_737
timestamp 1626908933
transform 1 0 24500 0 1 8658
box -100 -49 100 49
use M1M2_PR  M1M2_PR_84
timestamp 1626908933
transform 1 0 24144 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_881
timestamp 1626908933
transform 1 0 24240 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2051
timestamp 1626908933
transform 1 0 24144 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2848
timestamp 1626908933
transform 1 0 24240 0 1 8917
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_223
timestamp 1626908933
transform 1 0 23904 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_945
timestamp 1626908933
transform 1 0 23904 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_48
timestamp 1626908933
transform -1 0 25440 0 -1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_9
timestamp 1626908933
transform -1 0 25440 0 -1 9324
box -38 -49 614 715
use M1M2_PR  M1M2_PR_2847
timestamp 1626908933
transform 1 0 24720 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2846
timestamp 1626908933
transform 1 0 24720 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_880
timestamp 1626908933
transform 1 0 24720 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_879
timestamp 1626908933
transform 1 0 24720 0 1 8769
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_841
timestamp 1626908933
transform 1 0 24672 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_240
timestamp 1626908933
transform 1 0 24672 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_961
timestamp 1626908933
transform 1 0 25680 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2928
timestamp 1626908933
transform 1 0 25680 0 1 8547
box -32 -32 32 32
use L1M1_PR  L1M1_PR_927
timestamp 1626908933
transform 1 0 25008 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2862
timestamp 1626908933
transform 1 0 25008 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_960
timestamp 1626908933
transform 1 0 25680 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_965
timestamp 1626908933
transform 1 0 25488 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2927
timestamp 1626908933
transform 1 0 25680 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2932
timestamp 1626908933
transform 1 0 25488 0 1 8917
box -32 -32 32 32
use L1M1_PR  L1M1_PR_929
timestamp 1626908933
transform 1 0 25200 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2864
timestamp 1626908933
transform 1 0 25200 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_118
timestamp 1626908933
transform 1 0 25440 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_716
timestamp 1626908933
transform 1 0 25440 0 -1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_195
timestamp 1626908933
transform 1 0 25968 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1024
timestamp 1626908933
transform 1 0 25776 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2130
timestamp 1626908933
transform 1 0 25968 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2959
timestamp 1626908933
transform 1 0 25776 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_959
timestamp 1626908933
transform 1 0 26256 0 1 9139
box -32 -32 32 32
use M1M2_PR  M1M2_PR_962
timestamp 1626908933
transform 1 0 26448 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2926
timestamp 1626908933
transform 1 0 26256 0 1 9139
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2929
timestamp 1626908933
transform 1 0 26448 0 1 8917
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_171
timestamp 1626908933
transform 1 0 25824 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_893
timestamp 1626908933
transform 1 0 25824 0 -1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2956
timestamp 1626908933
transform 1 0 26736 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1021
timestamp 1626908933
transform 1 0 26736 0 1 9065
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2145
timestamp 1626908933
transform 1 0 26736 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2144
timestamp 1626908933
transform 1 0 26736 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_178
timestamp 1626908933
transform 1 0 26736 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_177
timestamp 1626908933
transform 1 0 26736 0 1 8769
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1752
timestamp 1626908933
transform 1 0 26592 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_761
timestamp 1626908933
transform 1 0 26592 0 -1 9324
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_713
timestamp 1626908933
transform 1 0 26900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_65
timestamp 1626908933
transform 1 0 26900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_713
timestamp 1626908933
transform 1 0 26900 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_65
timestamp 1626908933
transform 1 0 26900 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2961
timestamp 1626908933
transform 1 0 26832 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1026
timestamp 1626908933
transform 1 0 26832 0 1 8917
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_86
timestamp 1626908933
transform 1 0 26688 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_25
timestamp 1626908933
transform 1 0 26688 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_762
timestamp 1626908933
transform 1 0 27360 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1753
timestamp 1626908933
transform 1 0 27360 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_194
timestamp 1626908933
transform 1 0 27024 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2129
timestamp 1626908933
transform 1 0 27024 0 1 8769
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_21
timestamp 1626908933
transform 1 0 26976 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_73
timestamp 1626908933
transform 1 0 26976 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_840
timestamp 1626908933
transform 1 0 27552 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_239
timestamp 1626908933
transform 1 0 27552 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_610
timestamp 1626908933
transform 1 0 27456 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_253
timestamp 1626908933
transform 1 0 27456 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2127
timestamp 1626908933
transform 1 0 28368 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_192
timestamp 1626908933
transform 1 0 28368 0 1 8399
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2845
timestamp 1626908933
transform 1 0 27792 0 1 8843
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2841
timestamp 1626908933
transform 1 0 28272 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_878
timestamp 1626908933
transform 1 0 27792 0 1 8843
box -32 -32 32 32
use M1M2_PR  M1M2_PR_874
timestamp 1626908933
transform 1 0 28272 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_851
timestamp 1626908933
transform 1 0 27744 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_129
timestamp 1626908933
transform 1 0 27744 0 -1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2860
timestamp 1626908933
transform 1 0 28656 0 1 8843
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2854
timestamp 1626908933
transform 1 0 28656 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_925
timestamp 1626908933
transform 1 0 28656 0 1 8843
box -29 -23 29 23
use L1M1_PR  L1M1_PR_919
timestamp 1626908933
transform 1 0 28656 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1754
timestamp 1626908933
transform 1 0 28512 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_763
timestamp 1626908933
transform 1 0 28512 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2858
timestamp 1626908933
transform 1 0 28848 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_923
timestamp 1626908933
transform 1 0 28848 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1451
timestamp 1626908933
transform 1 0 28896 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_460
timestamp 1626908933
transform 1 0 28896 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_80
timestamp 1626908933
transform -1 0 28896 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_18
timestamp 1626908933
transform -1 0 28896 0 -1 9324
box -38 -49 326 715
use M1M2_PR  M1M2_PR_876
timestamp 1626908933
transform 1 0 28944 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2843
timestamp 1626908933
transform 1 0 28944 0 1 8991
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_41
timestamp 1626908933
transform 1 0 29300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_689
timestamp 1626908933
transform 1 0 29300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_41
timestamp 1626908933
transform 1 0 29300 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_689
timestamp 1626908933
transform 1 0 29300 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_94
timestamp 1626908933
transform 1 0 28992 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_816
timestamp 1626908933
transform 1 0 28992 0 -1 9324
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3755
timestamp 1626908933
transform 1 0 29616 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1788
timestamp 1626908933
transform 1 0 29616 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_839
timestamp 1626908933
transform 1 0 29760 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_238
timestamp 1626908933
transform 1 0 29760 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_630
timestamp 1626908933
transform 1 0 29952 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_32
timestamp 1626908933
transform 1 0 29952 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_777
timestamp 1626908933
transform 1 0 30336 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_55
timestamp 1626908933
transform 1 0 30336 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_608
timestamp 1626908933
transform 1 0 31104 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_10
timestamp 1626908933
transform 1 0 31104 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_459
timestamp 1626908933
transform 1 0 31488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1450
timestamp 1626908933
transform 1 0 31488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_252
timestamp 1626908933
transform 1 0 31680 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_609
timestamp 1626908933
transform 1 0 31680 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_764
timestamp 1626908933
transform 1 0 31584 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1755
timestamp 1626908933
transform 1 0 31584 0 -1 9324
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_17
timestamp 1626908933
transform 1 0 31700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_665
timestamp 1626908933
transform 1 0 31700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_17
timestamp 1626908933
transform 1 0 31700 0 1 8658
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_665
timestamp 1626908933
transform 1 0 31700 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_423
timestamp 1626908933
transform 1 0 31776 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1024
timestamp 1626908933
transform 1 0 31776 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3753
timestamp 1626908933
transform 1 0 31824 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1786
timestamp 1626908933
transform 1 0 31824 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1756
timestamp 1626908933
transform 1 0 31968 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_765
timestamp 1626908933
transform 1 0 31968 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_251
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_608
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_237
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_424
timestamp 1626908933
transform 1 0 0 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_838
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1025
timestamp 1626908933
transform 1 0 0 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_766
timestamp 1626908933
transform 1 0 192 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1757
timestamp 1626908933
transform 1 0 192 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_695
timestamp 1626908933
transform 1 0 576 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1417
timestamp 1626908933
transform 1 0 576 0 1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1771
timestamp 1626908933
transform 1 0 1104 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3706
timestamp 1626908933
transform 1 0 1104 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3221
timestamp 1626908933
transform 1 0 1488 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1286
timestamp 1626908933
transform 1 0 1488 0 1 9435
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3181
timestamp 1626908933
transform 1 0 1488 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1214
timestamp 1626908933
transform 1 0 1488 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3142
timestamp 1626908933
transform 1 0 1392 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1207
timestamp 1626908933
transform 1 0 1392 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3104
timestamp 1626908933
transform 1 0 1488 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1137
timestamp 1626908933
transform 1 0 1488 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_118
timestamp 1626908933
transform 1 0 1344 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_56
timestamp 1626908933
transform 1 0 1344 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_767
timestamp 1626908933
transform 1 0 1632 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1758
timestamp 1626908933
transform 1 0 1632 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_336
timestamp 1626908933
transform 1 0 1680 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2271
timestamp 1626908933
transform 1 0 1680 0 1 9435
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_641
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1289
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_641
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1289
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3727
timestamp 1626908933
transform 1 0 1872 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1760
timestamp 1626908933
transform 1 0 1872 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3714
timestamp 1626908933
transform 1 0 2064 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1779
timestamp 1626908933
transform 1 0 2064 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3731
timestamp 1626908933
transform 1 0 2064 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1764
timestamp 1626908933
transform 1 0 2064 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3700
timestamp 1626908933
transform 1 0 1776 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1765
timestamp 1626908933
transform 1 0 1776 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3705
timestamp 1626908933
transform 1 0 1968 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1770
timestamp 1626908933
transform 1 0 1968 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3726
timestamp 1626908933
transform 1 0 1872 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1759
timestamp 1626908933
transform 1 0 1872 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3730
timestamp 1626908933
transform 1 0 2064 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1763
timestamp 1626908933
transform 1 0 2064 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3708
timestamp 1626908933
transform 1 0 2352 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1773
timestamp 1626908933
transform 1 0 2352 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2277
timestamp 1626908933
transform 1 0 2256 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_310
timestamp 1626908933
transform 1 0 2256 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3699
timestamp 1626908933
transform 1 0 2352 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3331
timestamp 1626908933
transform 1 0 2160 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1764
timestamp 1626908933
transform 1 0 2352 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1396
timestamp 1626908933
transform 1 0 2160 0 1 9879
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3721
timestamp 1626908933
transform 1 0 2448 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1754
timestamp 1626908933
transform 1 0 2448 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1026
timestamp 1626908933
transform 1 0 2208 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_425
timestamp 1626908933
transform 1 0 2208 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_2
timestamp 1626908933
transform 1 0 2400 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_5
timestamp 1626908933
transform 1 0 2400 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_23
timestamp 1626908933
transform 1 0 1728 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_48
timestamp 1626908933
transform 1 0 1728 0 1 9324
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3713
timestamp 1626908933
transform 1 0 2544 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3338
timestamp 1626908933
transform 1 0 2736 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1778
timestamp 1626908933
transform 1 0 2544 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1403
timestamp 1626908933
transform 1 0 2736 0 1 9731
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_458
timestamp 1626908933
transform 1 0 2880 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1449
timestamp 1626908933
transform 1 0 2880 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1761
timestamp 1626908933
transform 1 0 3312 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1762
timestamp 1626908933
transform 1 0 3312 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3728
timestamp 1626908933
transform 1 0 3312 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3729
timestamp 1626908933
transform 1 0 3312 0 1 9213
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1265
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_617
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1265
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_617
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1599
timestamp 1626908933
transform 1 0 3504 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3566
timestamp 1626908933
transform 1 0 3504 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1152
timestamp 1626908933
transform 1 0 3792 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3119
timestamp 1626908933
transform 1 0 3792 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1223
timestamp 1626908933
transform 1 0 3792 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3158
timestamp 1626908933
transform 1 0 3792 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1692
timestamp 1626908933
transform 1 0 3984 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3627
timestamp 1626908933
transform 1 0 3984 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1316
timestamp 1626908933
transform 1 0 3888 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3283
timestamp 1626908933
transform 1 0 3888 0 1 9879
box -32 -32 32 32
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_7
timestamp 1626908933
transform 1 0 3744 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_2
timestamp 1626908933
transform 1 0 3744 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_647
timestamp 1626908933
transform 1 0 2976 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1369
timestamp 1626908933
transform 1 0 2976 0 1 9324
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1331
timestamp 1626908933
transform 1 0 4560 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3298
timestamp 1626908933
transform 1 0 4560 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1772
timestamp 1626908933
transform 1 0 4176 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3707
timestamp 1626908933
transform 1 0 4176 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3340
timestamp 1626908933
transform 1 0 5040 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1405
timestamp 1626908933
transform 1 0 5040 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3291
timestamp 1626908933
transform 1 0 5136 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3289
timestamp 1626908933
transform 1 0 4944 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1324
timestamp 1626908933
transform 1 0 5136 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1322
timestamp 1626908933
transform 1 0 4944 0 1 9731
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_607
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_250
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2069
timestamp 1626908933
transform 1 0 5520 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_134
timestamp 1626908933
transform 1 0 5520 0 1 9435
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1103
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_505
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_622
timestamp 1626908933
transform 1 0 4224 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1344
timestamp 1626908933
transform 1 0 4224 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_26
timestamp 1626908933
transform -1 0 7680 0 1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_1
timestamp 1626908933
transform -1 0 7680 0 1 9324
box -38 -49 2246 715
use M1M2_PR  M1M2_PR_1320
timestamp 1626908933
transform 1 0 5808 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3287
timestamp 1626908933
transform 1 0 5808 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1400
timestamp 1626908933
transform 1 0 6192 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3335
timestamp 1626908933
transform 1 0 6192 0 1 9213
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_593
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1241
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_593
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1241
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_121
timestamp 1626908933
transform 1 0 6864 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2088
timestamp 1626908933
transform 1 0 6864 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1616
timestamp 1626908933
transform 1 0 7440 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3551
timestamp 1626908933
transform 1 0 7440 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1529
timestamp 1626908933
transform 1 0 7632 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3496
timestamp 1626908933
transform 1 0 7632 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1479
timestamp 1626908933
transform 1 0 8016 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3446
timestamp 1626908933
transform 1 0 8016 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1565
timestamp 1626908933
transform 1 0 8112 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3500
timestamp 1626908933
transform 1 0 8112 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1944
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3911
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1913
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3848
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1528
timestamp 1626908933
transform 1 0 7632 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3495
timestamp 1626908933
transform 1 0 7632 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1566
timestamp 1626908933
transform 1 0 7728 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1615
timestamp 1626908933
transform 1 0 7632 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3501
timestamp 1626908933
transform 1 0 7728 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3550
timestamp 1626908933
transform 1 0 7632 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1478
timestamp 1626908933
transform 1 0 8016 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3445
timestamp 1626908933
transform 1 0 8016 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1671
timestamp 1626908933
transform 1 0 8208 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3638
timestamp 1626908933
transform 1 0 8208 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1756
timestamp 1626908933
transform 1 0 8112 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3691
timestamp 1626908933
transform 1 0 8112 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_25
timestamp 1626908933
transform 1 0 7680 0 1 9324
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_1
timestamp 1626908933
transform 1 0 7680 0 1 9324
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1217
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_569
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1217
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_569
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3701
timestamp 1626908933
transform 1 0 8400 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1988
timestamp 1626908933
transform 1 0 9072 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1734
timestamp 1626908933
transform 1 0 8400 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_21
timestamp 1626908933
transform 1 0 9072 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1957
timestamp 1626908933
transform 1 0 9936 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_22
timestamp 1626908933
transform 1 0 9936 0 1 9435
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2600
timestamp 1626908933
transform 1 0 9456 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_633
timestamp 1626908933
transform 1 0 9456 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_606
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_249
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1984
timestamp 1626908933
transform 1 0 10608 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_17
timestamp 1626908933
transform 1 0 10608 0 1 9435
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1023
timestamp 1626908933
transform 1 0 10080 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_425
timestamp 1626908933
transform 1 0 10080 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1241
timestamp 1626908933
transform 1 0 10464 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_519
timestamp 1626908933
transform 1 0 10464 0 1 9324
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1193
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_545
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1193
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_545
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2896
timestamp 1626908933
transform 1 0 11184 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_929
timestamp 1626908933
transform 1 0 11184 0 1 9213
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1759
timestamp 1626908933
transform 1 0 11232 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_768
timestamp 1626908933
transform 1 0 11232 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2576
timestamp 1626908933
transform 1 0 11376 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_641
timestamp 1626908933
transform 1 0 11376 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2619
timestamp 1626908933
transform 1 0 11472 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_684
timestamp 1626908933
transform 1 0 11472 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2634
timestamp 1626908933
transform 1 0 11472 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_667
timestamp 1626908933
transform 1 0 11472 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_631
timestamp 1626908933
transform 1 0 11568 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_773
timestamp 1626908933
transform 1 0 11760 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2598
timestamp 1626908933
transform 1 0 11568 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2740
timestamp 1626908933
transform 1 0 11760 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_789
timestamp 1626908933
transform 1 0 11568 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_803
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2724
timestamp 1626908933
transform 1 0 11568 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2738
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_486
timestamp 1626908933
transform 1 0 11712 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1208
timestamp 1626908933
transform 1 0 11712 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_5
timestamp 1626908933
transform -1 0 11712 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_13
timestamp 1626908933
transform -1 0 11712 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nand4_1  sky130_fd_sc_hs__nand4_1_5
timestamp 1626908933
transform -1 0 13152 0 1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__nand4_1  sky130_fd_sc_hs__nand4_1_2
timestamp 1626908933
transform -1 0 13152 0 1 9324
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2723
timestamp 1626908933
transform 1 0 12720 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2722
timestamp 1626908933
transform 1 0 12528 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_788
timestamp 1626908933
transform 1 0 12720 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_787
timestamp 1626908933
transform 1 0 12528 0 1 9879
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1760
timestamp 1626908933
transform 1 0 12480 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_769
timestamp 1626908933
transform 1 0 12480 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2725
timestamp 1626908933
transform 1 0 12912 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_790
timestamp 1626908933
transform 1 0 12912 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2727
timestamp 1626908933
transform 1 0 12816 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_760
timestamp 1626908933
transform 1 0 12816 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2569
timestamp 1626908933
transform 1 0 13008 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_634
timestamp 1626908933
transform 1 0 13008 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2591
timestamp 1626908933
transform 1 0 13008 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_624
timestamp 1626908933
transform 1 0 13008 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2648
timestamp 1626908933
transform 1 0 13104 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_713
timestamp 1626908933
transform 1 0 13104 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_457
timestamp 1626908933
transform 1 0 13536 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1448
timestamp 1626908933
transform 1 0 13536 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_353
timestamp 1626908933
transform 1 0 13152 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_951
timestamp 1626908933
transform 1 0 13152 0 1 9324
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1169
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_521
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1169
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_521
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1167
timestamp 1626908933
transform 1 0 13632 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_445
timestamp 1626908933
transform 1 0 13632 0 1 9324
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1515
timestamp 1626908933
transform 1 0 13968 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3482
timestamp 1626908933
transform 1 0 13968 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_983
timestamp 1626908933
transform 1 0 13872 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1601
timestamp 1626908933
transform 1 0 14160 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2918
timestamp 1626908933
transform 1 0 13872 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3536
timestamp 1626908933
transform 1 0 14160 0 1 9213
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_236
timestamp 1626908933
transform 1 0 14400 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_837
timestamp 1626908933
transform 1 0 14400 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_334
timestamp 1626908933
transform 1 0 14592 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_932
timestamp 1626908933
transform 1 0 14592 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1447
timestamp 1626908933
transform 1 0 15456 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_456
timestamp 1626908933
transform 1 0 15456 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_921
timestamp 1626908933
transform 1 0 15072 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_323
timestamp 1626908933
transform 1 0 15072 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_605
timestamp 1626908933
transform 1 0 14976 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_248
timestamp 1626908933
transform 1 0 14976 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_14
timestamp 1626908933
transform 1 0 15600 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1981
timestamp 1626908933
transform 1 0 15600 0 1 9435
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_455
timestamp 1626908933
transform 1 0 16320 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1446
timestamp 1626908933
transform 1 0 16320 0 1 9324
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_497
timestamp 1626908933
transform 1 0 16100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1145
timestamp 1626908933
transform 1 0 16100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_497
timestamp 1626908933
transform 1 0 16100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1145
timestamp 1626908933
transform 1 0 16100 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_411
timestamp 1626908933
transform 1 0 15552 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1133
timestamp 1626908933
transform 1 0 15552 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_895
timestamp 1626908933
transform 1 0 16416 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_297
timestamp 1626908933
transform 1 0 16416 0 1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2675
timestamp 1626908933
transform 1 0 17328 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2662
timestamp 1626908933
transform 1 0 16848 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_708
timestamp 1626908933
transform 1 0 17328 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_695
timestamp 1626908933
transform 1 0 16848 0 1 9435
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1104
timestamp 1626908933
transform 1 0 16800 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_382
timestamp 1626908933
transform 1 0 16800 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_235
timestamp 1626908933
transform 1 0 17568 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_426
timestamp 1626908933
transform 1 0 17760 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_836
timestamp 1626908933
transform 1 0 17568 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1027
timestamp 1626908933
transform 1 0 17760 0 1 9324
box -38 -49 230 715
use L1M1_PR  L1M1_PR_2649
timestamp 1626908933
transform 1 0 18000 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_714
timestamp 1626908933
transform 1 0 18000 0 1 9435
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1761
timestamp 1626908933
transform 1 0 17952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_770
timestamp 1626908933
transform 1 0 17952 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2647
timestamp 1626908933
transform 1 0 18192 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2646
timestamp 1626908933
transform 1 0 18096 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_712
timestamp 1626908933
transform 1 0 18192 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_711
timestamp 1626908933
transform 1 0 18096 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2726
timestamp 1626908933
transform 1 0 18192 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_759
timestamp 1626908933
transform 1 0 18192 0 1 9879
box -32 -32 32 32
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_1
timestamp 1626908933
transform -1 0 18432 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_9
timestamp 1626908933
transform -1 0 18432 0 1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_694
timestamp 1626908933
transform 1 0 18288 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2661
timestamp 1626908933
transform 1 0 18288 0 1 9213
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_473
timestamp 1626908933
transform 1 0 18500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1121
timestamp 1626908933
transform 1 0 18500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_473
timestamp 1626908933
transform 1 0 18500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1121
timestamp 1626908933
transform 1 0 18500 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_693
timestamp 1626908933
transform 1 0 18288 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2660
timestamp 1626908933
transform 1 0 18288 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_421
timestamp 1626908933
transform 1 0 18288 0 1 9805
box -29 -23 29 23
use L1M1_PR  L1M1_PR_710
timestamp 1626908933
transform 1 0 18384 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2356
timestamp 1626908933
transform 1 0 18288 0 1 9805
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2645
timestamp 1626908933
transform 1 0 18384 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_454
timestamp 1626908933
transform 1 0 18432 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1445
timestamp 1626908933
transform 1 0 18432 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_597
timestamp 1626908933
transform 1 0 18960 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2564
timestamp 1626908933
transform 1 0 18960 0 1 9509
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_337
timestamp 1626908933
transform 1 0 18528 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1059
timestamp 1626908933
transform 1 0 18528 0 1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2461
timestamp 1626908933
transform 1 0 19248 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_526
timestamp 1626908933
transform 1 0 19248 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2145
timestamp 1626908933
transform 1 0 19344 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_210
timestamp 1626908933
transform 1 0 19344 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2496
timestamp 1626908933
transform 1 0 19344 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2158
timestamp 1626908933
transform 1 0 19248 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_529
timestamp 1626908933
transform 1 0 19344 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_191
timestamp 1626908933
transform 1 0 19248 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_76
timestamp 1626908933
transform 1 0 19296 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_14
timestamp 1626908933
transform 1 0 19296 0 1 9324
box -38 -49 326 715
use M1M2_PR  M1M2_PR_425
timestamp 1626908933
transform 1 0 19536 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_733
timestamp 1626908933
transform 1 0 19536 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2392
timestamp 1626908933
transform 1 0 19536 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2700
timestamp 1626908933
transform 1 0 19536 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_528
timestamp 1626908933
transform 1 0 19440 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_756
timestamp 1626908933
transform 1 0 19536 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2463
timestamp 1626908933
transform 1 0 19440 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2691
timestamp 1626908933
transform 1 0 19536 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_247
timestamp 1626908933
transform 1 0 19968 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_604
timestamp 1626908933
transform 1 0 19968 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_427
timestamp 1626908933
transform 1 0 20064 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1028
timestamp 1626908933
transform 1 0 20064 0 1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_526
timestamp 1626908933
transform 1 0 20112 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_527
timestamp 1626908933
transform 1 0 20112 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2493
timestamp 1626908933
transform 1 0 20112 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2494
timestamp 1626908933
transform 1 0 20112 0 1 9213
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_221
timestamp 1626908933
transform 1 0 19584 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_819
timestamp 1626908933
transform 1 0 19584 0 1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2460
timestamp 1626908933
transform 1 0 20208 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_525
timestamp 1626908933
transform 1 0 20208 0 1 9435
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2390
timestamp 1626908933
transform 1 0 20304 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_423
timestamp 1626908933
transform 1 0 20304 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2353
timestamp 1626908933
transform 1 0 20400 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_418
timestamp 1626908933
transform 1 0 20400 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2458
timestamp 1626908933
transform 1 0 20496 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_523
timestamp 1626908933
transform 1 0 20496 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2456
timestamp 1626908933
transform 1 0 20592 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_521
timestamp 1626908933
transform 1 0 20592 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2492
timestamp 1626908933
transform 1 0 20496 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_525
timestamp 1626908933
transform 1 0 20496 0 1 9657
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1097
timestamp 1626908933
transform 1 0 20900 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_449
timestamp 1626908933
transform 1 0 20900 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1097
timestamp 1626908933
transform 1 0 20900 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_449
timestamp 1626908933
transform 1 0 20900 0 1 9324
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2462
timestamp 1626908933
transform 1 0 20880 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_527
timestamp 1626908933
transform 1 0 20880 0 1 9879
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2489
timestamp 1626908933
transform 1 0 20688 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_522
timestamp 1626908933
transform 1 0 20688 0 1 9583
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_835
timestamp 1626908933
transform 1 0 20832 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_234
timestamp 1626908933
transform 1 0 20832 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_285
timestamp 1626908933
transform 1 0 21024 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1007
timestamp 1626908933
transform 1 0 21024 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__a31oi_1  sky130_fd_sc_hs__a31oi_1_0
timestamp 1626908933
transform 1 0 20256 0 1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__a31oi_1  sky130_fd_sc_hs__a31oi_1_1
timestamp 1626908933
transform 1 0 20256 0 1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__nand4_1  sky130_fd_sc_hs__nand4_1_4
timestamp 1626908933
transform 1 0 21792 0 1 9324
box -38 -49 614 715
use sky130_fd_sc_hs__nand4_1  sky130_fd_sc_hs__nand4_1_1
timestamp 1626908933
transform 1 0 21792 0 1 9324
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2665
timestamp 1626908933
transform 1 0 21744 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2043
timestamp 1626908933
transform 1 0 21072 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_730
timestamp 1626908933
transform 1 0 21744 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_108
timestamp 1626908933
transform 1 0 21072 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2061
timestamp 1626908933
transform 1 0 21456 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_94
timestamp 1626908933
transform 1 0 21456 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2541
timestamp 1626908933
transform 1 0 22032 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2506
timestamp 1626908933
transform 1 0 21936 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_606
timestamp 1626908933
transform 1 0 22032 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_571
timestamp 1626908933
transform 1 0 21936 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2041
timestamp 1626908933
transform 1 0 22224 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_106
timestamp 1626908933
transform 1 0 22224 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_713
timestamp 1626908933
transform 1 0 22224 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2680
timestamp 1626908933
transform 1 0 22224 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_735
timestamp 1626908933
transform 1 0 22224 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2670
timestamp 1626908933
transform 1 0 22224 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_711
timestamp 1626908933
transform 1 0 22320 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2678
timestamp 1626908933
transform 1 0 22320 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_732
timestamp 1626908933
transform 1 0 22320 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2667
timestamp 1626908933
transform 1 0 22320 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_549
timestamp 1626908933
transform 1 0 22512 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2516
timestamp 1626908933
transform 1 0 22512 0 1 9731
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_834
timestamp 1626908933
transform 1 0 22368 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_233
timestamp 1626908933
transform 1 0 22368 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_253
timestamp 1626908933
transform 1 0 22560 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_975
timestamp 1626908933
transform 1 0 22560 0 1 9324
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1073
timestamp 1626908933
transform 1 0 23300 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_425
timestamp 1626908933
transform 1 0 23300 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1073
timestamp 1626908933
transform 1 0 23300 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_425
timestamp 1626908933
transform 1 0 23300 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2510
timestamp 1626908933
transform 1 0 23088 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_543
timestamp 1626908933
transform 1 0 23088 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2535
timestamp 1626908933
transform 1 0 23280 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_568
timestamp 1626908933
transform 1 0 23280 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_833
timestamp 1626908933
transform 1 0 23328 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_232
timestamp 1626908933
transform 1 0 23328 0 1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_551
timestamp 1626908933
transform 1 0 23664 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2518
timestamp 1626908933
transform 1 0 23664 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_545
timestamp 1626908933
transform 1 0 23664 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_553
timestamp 1626908933
transform 1 0 23760 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_558
timestamp 1626908933
transform 1 0 23472 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2480
timestamp 1626908933
transform 1 0 23664 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2488
timestamp 1626908933
transform 1 0 23760 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2493
timestamp 1626908933
transform 1 0 23472 0 1 9879
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_2
timestamp 1626908933
transform -1 0 23904 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_64
timestamp 1626908933
transform -1 0 23904 0 1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2491
timestamp 1626908933
transform 1 0 23856 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_556
timestamp 1626908933
transform 1 0 23856 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2520
timestamp 1626908933
transform 1 0 23856 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_553
timestamp 1626908933
transform 1 0 23856 0 1 9879
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_944
timestamp 1626908933
transform 1 0 23904 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_222
timestamp 1626908933
transform 1 0 23904 0 1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2039
timestamp 1626908933
transform 1 0 24816 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_104
timestamp 1626908933
transform 1 0 24816 0 1 9213
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1762
timestamp 1626908933
transform 1 0 24864 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_771
timestamp 1626908933
transform 1 0 24864 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1029
timestamp 1626908933
transform 1 0 24672 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_428
timestamp 1626908933
transform 1 0 24672 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_246
timestamp 1626908933
transform 1 0 24960 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_603
timestamp 1626908933
transform 1 0 24960 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_92
timestamp 1626908933
transform 1 0 25104 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_93
timestamp 1626908933
transform 1 0 25104 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2059
timestamp 1626908933
transform 1 0 25104 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2060
timestamp 1626908933
transform 1 0 25104 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_103
timestamp 1626908933
transform 1 0 25104 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2038
timestamp 1626908933
transform 1 0 25104 0 1 9435
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1444
timestamp 1626908933
transform 1 0 25392 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1445
timestamp 1626908933
transform 1 0 25392 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3411
timestamp 1626908933
transform 1 0 25392 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3412
timestamp 1626908933
transform 1 0 25392 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1530
timestamp 1626908933
transform 1 0 25392 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3465
timestamp 1626908933
transform 1 0 25392 0 1 9213
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_401
timestamp 1626908933
transform 1 0 25700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1049
timestamp 1626908933
transform 1 0 25700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_401
timestamp 1626908933
transform 1 0 25700 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1049
timestamp 1626908933
transform 1 0 25700 0 1 9324
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3670
timestamp 1626908933
transform 1 0 26928 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3464
timestamp 1626908933
transform 1 0 27312 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1735
timestamp 1626908933
transform 1 0 26928 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1529
timestamp 1626908933
transform 1 0 27312 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3620
timestamp 1626908933
transform 1 0 27408 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1653
timestamp 1626908933
transform 1 0 27408 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_685
timestamp 1626908933
transform 1 0 27360 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_87
timestamp 1626908933
transform 1 0 27360 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_42
timestamp 1626908933
transform -1 0 27360 0 1 9324
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_18
timestamp 1626908933
transform -1 0 27360 0 1 9324
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1025
timestamp 1626908933
transform 1 0 28100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_377
timestamp 1626908933
transform 1 0 28100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1025
timestamp 1626908933
transform 1 0 28100 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_377
timestamp 1626908933
transform 1 0 28100 0 1 9324
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2861
timestamp 1626908933
transform 1 0 27792 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_926
timestamp 1626908933
transform 1 0 27792 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2844
timestamp 1626908933
transform 1 0 27792 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_877
timestamp 1626908933
transform 1 0 27792 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2859
timestamp 1626908933
transform 1 0 27984 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_924
timestamp 1626908933
transform 1 0 27984 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3466
timestamp 1626908933
transform 1 0 27792 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1531
timestamp 1626908933
transform 1 0 27792 0 1 9879
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3414
timestamp 1626908933
transform 1 0 27696 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1447
timestamp 1626908933
transform 1 0 27696 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3646
timestamp 1626908933
transform 1 0 27888 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1679
timestamp 1626908933
transform 1 0 27888 0 1 9805
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_231
timestamp 1626908933
transform 1 0 28128 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_832
timestamp 1626908933
transform 1 0 28128 0 1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_873
timestamp 1626908933
transform 1 0 28272 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2840
timestamp 1626908933
transform 1 0 28272 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_921
timestamp 1626908933
transform 1 0 28080 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2856
timestamp 1626908933
transform 1 0 28080 0 1 9583
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_109
timestamp 1626908933
transform 1 0 28320 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_831
timestamp 1626908933
transform 1 0 28320 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_22
timestamp 1626908933
transform -1 0 28128 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_84
timestamp 1626908933
transform -1 0 28128 0 1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2857
timestamp 1626908933
transform 1 0 29232 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_922
timestamp 1626908933
transform 1 0 29232 0 1 9731
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2842
timestamp 1626908933
transform 1 0 28944 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_875
timestamp 1626908933
transform 1 0 28944 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_25
timestamp 1626908933
transform 1 0 29088 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_94
timestamp 1626908933
transform 1 0 29088 0 1 9324
box -38 -49 518 715
use M1M2_PR  M1M2_PR_89
timestamp 1626908933
transform 1 0 29520 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2056
timestamp 1626908933
transform 1 0 29520 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_100
timestamp 1626908933
transform 1 0 29424 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2035
timestamp 1626908933
transform 1 0 29424 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_245
timestamp 1626908933
transform 1 0 29952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_602
timestamp 1626908933
transform 1 0 29952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_230
timestamp 1626908933
transform 1 0 30048 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_831
timestamp 1626908933
transform 1 0 30048 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_45
timestamp 1626908933
transform 1 0 29568 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_643
timestamp 1626908933
transform 1 0 29568 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1444
timestamp 1626908933
transform 1 0 30240 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_453
timestamp 1626908933
transform 1 0 30240 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_776
timestamp 1626908933
transform 1 0 30336 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_54
timestamp 1626908933
transform 1 0 30336 0 1 9324
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1001
timestamp 1626908933
transform 1 0 30500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_353
timestamp 1626908933
transform 1 0 30500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1001
timestamp 1626908933
transform 1 0 30500 0 1 9324
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_353
timestamp 1626908933
transform 1 0 30500 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1443
timestamp 1626908933
transform 1 0 31104 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_452
timestamp 1626908933
transform 1 0 31104 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_738
timestamp 1626908933
transform 1 0 31200 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_16
timestamp 1626908933
transform 1 0 31200 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1763
timestamp 1626908933
transform 1 0 31968 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_772
timestamp 1626908933
transform 1 0 31968 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1773
timestamp 1626908933
transform 1 0 192 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_782
timestamp 1626908933
transform 1 0 192 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1427
timestamp 1626908933
transform 1 0 384 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_436
timestamp 1626908933
transform 1 0 384 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_594
timestamp 1626908933
transform 1 0 288 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_237
timestamp 1626908933
transform 1 0 288 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1037
timestamp 1626908933
transform 1 0 0 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_830
timestamp 1626908933
transform 1 0 0 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_436
timestamp 1626908933
transform 1 0 0 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_229
timestamp 1626908933
transform 1 0 0 0 -1 10656
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_328
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_976
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_328
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_976
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_715
timestamp 1626908933
transform 1 0 192 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1437
timestamp 1626908933
transform 1 0 192 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_592
timestamp 1626908933
transform 1 0 480 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1190
timestamp 1626908933
transform 1 0 480 0 1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3885
timestamp 1626908933
transform 1 0 1008 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1918
timestamp 1626908933
transform 1 0 1008 0 1 10249
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1774
timestamp 1626908933
transform 1 0 960 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1426
timestamp 1626908933
transform 1 0 864 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_783
timestamp 1626908933
transform 1 0 960 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_435
timestamp 1626908933
transform 1 0 864 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3702
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1767
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3735
timestamp 1626908933
transform 1 0 1104 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3722
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1768
timestamp 1626908933
transform 1 0 1104 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1755
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_121
timestamp 1626908933
transform 1 0 1056 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_59
timestamp 1626908933
transform 1 0 1056 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_829
timestamp 1626908933
transform 1 0 960 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_228
timestamp 1626908933
transform 1 0 960 0 -1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3717
timestamp 1626908933
transform 1 0 1392 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1782
timestamp 1626908933
transform 1 0 1392 0 1 10545
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1425
timestamp 1626908933
transform 1 0 1344 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_434
timestamp 1626908933
transform 1 0 1344 0 1 10656
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1288
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_640
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1288
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_640
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3823
timestamp 1626908933
transform 1 0 1584 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1888
timestamp 1626908933
transform 1 0 1584 0 1 10249
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3103
timestamp 1626908933
transform 1 0 1488 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1136
timestamp 1626908933
transform 1 0 1488 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3141
timestamp 1626908933
transform 1 0 1680 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1206
timestamp 1626908933
transform 1 0 1680 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_682
timestamp 1626908933
transform 1 0 1440 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1404
timestamp 1626908933
transform 1 0 1440 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__or3b_2  sky130_fd_sc_hs__or3b_2_0
timestamp 1626908933
transform 1 0 1152 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__or3b_2  sky130_fd_sc_hs__or3b_2_1
timestamp 1626908933
transform 1 0 1152 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_451
timestamp 1626908933
transform 1 0 1920 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1442
timestamp 1626908933
transform 1 0 1920 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1424
timestamp 1626908933
transform 1 0 2208 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_433
timestamp 1626908933
transform 1 0 2208 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3720
timestamp 1626908933
transform 1 0 2448 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3302
timestamp 1626908933
transform 1 0 2448 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1753
timestamp 1626908933
transform 1 0 2448 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1335
timestamp 1626908933
transform 1 0 2448 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1441
timestamp 1626908933
transform 1 0 2400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_450
timestamp 1626908933
transform 1 0 2400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_601
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_244
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_656
timestamp 1626908933
transform 1 0 2304 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1378
timestamp 1626908933
transform 1 0 2304 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_555
timestamp 1626908933
transform 1 0 2016 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1153
timestamp 1626908933
transform 1 0 2016 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1030
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_429
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_952
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_304
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_952
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_304
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3698
timestamp 1626908933
transform 1 0 2928 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3348
timestamp 1626908933
transform 1 0 2832 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1763
timestamp 1626908933
transform 1 0 2928 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1413
timestamp 1626908933
transform 1 0 2832 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3884
timestamp 1626908933
transform 1 0 3216 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3718
timestamp 1626908933
transform 1 0 3120 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1917
timestamp 1626908933
transform 1 0 3216 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1751
timestamp 1626908933
transform 1 0 3120 0 1 10101
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1440
timestamp 1626908933
transform 1 0 3264 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_449
timestamp 1626908933
transform 1 0 3264 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_68
timestamp 1626908933
transform 1 0 2784 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_137
timestamp 1626908933
transform 1 0 2784 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_448
timestamp 1626908933
transform 1 0 4128 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1439
timestamp 1626908933
transform 1 0 4128 0 -1 10656
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_616
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1264
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_616
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1264
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_646
timestamp 1626908933
transform 1 0 3360 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1368
timestamp 1626908933
transform 1 0 3360 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_524
timestamp 1626908933
transform 1 0 4224 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1122
timestamp 1626908933
transform 1 0 4224 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_227
timestamp 1626908933
transform 1 0 4608 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_437
timestamp 1626908933
transform 1 0 4800 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_828
timestamp 1626908933
transform 1 0 4608 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1038
timestamp 1626908933
transform 1 0 4800 0 1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1330
timestamp 1626908933
transform 1 0 4560 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3297
timestamp 1626908933
transform 1 0 4560 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3407
timestamp 1626908933
transform 1 0 4848 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1472
timestamp 1626908933
transform 1 0 4848 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3358
timestamp 1626908933
transform 1 0 4848 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1391
timestamp 1626908933
transform 1 0 4848 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_822
timestamp 1626908933
transform 1 0 5088 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_221
timestamp 1626908933
transform 1 0 5088 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_593
timestamp 1626908933
transform 1 0 4992 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_236
timestamp 1626908933
transform 1 0 4992 0 1 10656
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_928
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_280
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_928
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_280
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3339
timestamp 1626908933
transform 1 0 5232 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1404
timestamp 1626908933
transform 1 0 5232 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3290
timestamp 1626908933
transform 1 0 5136 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1323
timestamp 1626908933
transform 1 0 5136 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_605
timestamp 1626908933
transform 1 0 5280 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1327
timestamp 1626908933
transform 1 0 5280 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_11
timestamp 1626908933
transform -1 0 4800 0 1 10656
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_5
timestamp 1626908933
transform -1 0 4800 0 1 10656
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_5
timestamp 1626908933
transform 1 0 4800 0 -1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_0
timestamp 1626908933
transform 1 0 4800 0 -1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_493
timestamp 1626908933
transform 1 0 6048 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1091
timestamp 1626908933
transform 1 0 6048 0 1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_324
timestamp 1626908933
transform 1 0 5904 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2291
timestamp 1626908933
transform 1 0 5904 0 1 10101
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1240
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_592
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1240
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_592
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2285
timestamp 1626908933
transform 1 0 6384 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_350
timestamp 1626908933
transform 1 0 6384 0 1 10101
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1423
timestamp 1626908933
transform 1 0 6432 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_432
timestamp 1626908933
transform 1 0 6432 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1031
timestamp 1626908933
transform 1 0 6720 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_430
timestamp 1626908933
transform 1 0 6720 0 -1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_2674
timestamp 1626908933
transform 1 0 6864 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_707
timestamp 1626908933
transform 1 0 6864 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1764
timestamp 1626908933
transform 1 0 6912 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_773
timestamp 1626908933
transform 1 0 6912 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_577
timestamp 1626908933
transform 1 0 6528 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1299
timestamp 1626908933
transform 1 0 6528 0 1 10656
box -38 -49 806 715
use L1M1_PR  L1M1_PR_949
timestamp 1626908933
transform 1 0 7056 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2884
timestamp 1626908933
transform 1 0 7056 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_901
timestamp 1626908933
transform 1 0 7152 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2868
timestamp 1626908933
transform 1 0 7152 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_727
timestamp 1626908933
transform 1 0 7248 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2662
timestamp 1626908933
transform 1 0 7248 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_903
timestamp 1626908933
transform 1 0 7056 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2870
timestamp 1626908933
transform 1 0 7056 0 1 10545
box -32 -32 32 32
use L1M1_PR  L1M1_PR_950
timestamp 1626908933
transform 1 0 7152 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2885
timestamp 1626908933
transform 1 0 7152 0 1 10545
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1032
timestamp 1626908933
transform 1 0 7296 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_431
timestamp 1626908933
transform 1 0 7296 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_600
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_243
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_101
timestamp 1626908933
transform -1 0 7296 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_39
timestamp 1626908933
transform -1 0 7296 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1068
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_470
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_904
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_256
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_904
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_256
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3503
timestamp 1626908933
transform 1 0 8112 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1568
timestamp 1626908933
transform 1 0 8112 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3637
timestamp 1626908933
transform 1 0 8208 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1670
timestamp 1626908933
transform 1 0 8208 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1765
timestamp 1626908933
transform 1 0 7968 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_774
timestamp 1626908933
transform 1 0 7968 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_89
timestamp 1626908933
transform -1 0 8352 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_27
timestamp 1626908933
transform -1 0 8352 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_558
timestamp 1626908933
transform 1 0 7296 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1280
timestamp 1626908933
transform 1 0 7296 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_24
timestamp 1626908933
transform 1 0 8064 0 -1 10656
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_0
timestamp 1626908933
transform 1 0 8064 0 -1 10656
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_1481
timestamp 1626908933
transform 1 0 8688 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1733
timestamp 1626908933
transform 1 0 8400 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3448
timestamp 1626908933
transform 1 0 8688 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3700
timestamp 1626908933
transform 1 0 8400 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1754
timestamp 1626908933
transform 1 0 8496 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3689
timestamp 1626908933
transform 1 0 8496 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_438
timestamp 1626908933
transform 1 0 9120 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1039
timestamp 1626908933
transform 1 0 9120 0 1 10656
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_568
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1216
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_568
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1216
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_10
timestamp 1626908933
transform 1 0 8352 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_33
timestamp 1626908933
transform 1 0 8352 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_784
timestamp 1626908933
transform 1 0 9312 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1775
timestamp 1626908933
transform 1 0 9312 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_235
timestamp 1626908933
transform 1 0 9984 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_592
timestamp 1626908933
transform 1 0 9984 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_785
timestamp 1626908933
transform 1 0 9888 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1776
timestamp 1626908933
transform 1 0 9888 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_20
timestamp 1626908933
transform 1 0 9936 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1987
timestamp 1626908933
transform 1 0 9936 0 1 10545
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_85
timestamp 1626908933
transform -1 0 9888 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_16
timestamp 1626908933
transform -1 0 9888 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_447
timestamp 1626908933
transform 1 0 10368 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1438
timestamp 1626908933
transform 1 0 10368 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_19
timestamp 1626908933
transform 1 0 10320 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1954
timestamp 1626908933
transform 1 0 10320 0 1 10545
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_232
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_880
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_232
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_880
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use M1M2_PR  M1M2_PR_16
timestamp 1626908933
transform 1 0 10608 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1983
timestamp 1626908933
transform 1 0 10608 0 1 10101
box -32 -32 32 32
use L1M1_PR  L1M1_PR_18
timestamp 1626908933
transform 1 0 10416 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1953
timestamp 1626908933
transform 1 0 10416 0 1 10101
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_518
timestamp 1626908933
transform 1 0 10464 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1240
timestamp 1626908933
transform 1 0 10464 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_408
timestamp 1626908933
transform 1 0 10464 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_424
timestamp 1626908933
transform 1 0 10080 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1006
timestamp 1626908933
transform 1 0 10464 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1022
timestamp 1626908933
transform 1 0 10080 0 1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2094
timestamp 1626908933
transform 1 0 10992 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_159
timestamp 1626908933
transform 1 0 10992 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2112
timestamp 1626908933
transform 1 0 10896 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_145
timestamp 1626908933
transform 1 0 10896 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_7
timestamp 1626908933
transform -1 0 11328 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_76
timestamp 1626908933
transform -1 0 11328 0 -1 10656
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1192
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_544
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1192
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_544
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2736
timestamp 1626908933
transform 1 0 11184 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_801
timestamp 1626908933
transform 1 0 11184 0 1 10545
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2738
timestamp 1626908933
transform 1 0 11568 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_771
timestamp 1626908933
transform 1 0 11568 0 1 10545
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_72
timestamp 1626908933
transform -1 0 12000 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_10
timestamp 1626908933
transform -1 0 12000 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_29
timestamp 1626908933
transform -1 0 12096 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_4
timestamp 1626908933
transform -1 0 12096 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_995
timestamp 1626908933
transform 1 0 11328 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_994
timestamp 1626908933
transform 1 0 11232 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_397
timestamp 1626908933
transform 1 0 11328 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_396
timestamp 1626908933
transform 1 0 11232 0 1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_772
timestamp 1626908933
transform 1 0 11760 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2739
timestamp 1626908933
transform 1 0 11760 0 1 10101
box -32 -32 32 32
use L1M1_PR  L1M1_PR_673
timestamp 1626908933
transform 1 0 11760 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_802
timestamp 1626908933
transform 1 0 11760 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2608
timestamp 1626908933
transform 1 0 11760 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2737
timestamp 1626908933
transform 1 0 11760 0 1 10101
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_446
timestamp 1626908933
transform 1 0 12000 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1437
timestamp 1626908933
transform 1 0 12000 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_66
timestamp 1626908933
transform 1 0 12048 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2001
timestamp 1626908933
transform 1 0 12048 0 1 10249
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_856
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_208
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_856
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_208
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2625
timestamp 1626908933
transform 1 0 12336 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_658
timestamp 1626908933
transform 1 0 12336 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_978
timestamp 1626908933
transform 1 0 12096 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_380
timestamp 1626908933
transform 1 0 12096 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_11
timestamp 1626908933
transform 1 0 12096 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_34
timestamp 1626908933
transform 1 0 12096 0 1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2025
timestamp 1626908933
transform 1 0 12720 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_58
timestamp 1626908933
transform 1 0 12720 0 1 10249
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1766
timestamp 1626908933
transform 1 0 12768 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_775
timestamp 1626908933
transform 1 0 12768 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1033
timestamp 1626908933
transform 1 0 12576 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_432
timestamp 1626908933
transform 1 0 12576 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_599
timestamp 1626908933
transform 1 0 12480 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_242
timestamp 1626908933
transform 1 0 12480 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2607
timestamp 1626908933
transform 1 0 12912 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2535
timestamp 1626908933
transform 1 0 13104 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1998
timestamp 1626908933
transform 1 0 13008 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_672
timestamp 1626908933
transform 1 0 12912 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_600
timestamp 1626908933
transform 1 0 13104 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_63
timestamp 1626908933
transform 1 0 13008 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2558
timestamp 1626908933
transform 1 0 13008 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_591
timestamp 1626908933
transform 1 0 13008 0 1 10545
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_69
timestamp 1626908933
transform 1 0 12864 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_68
timestamp 1626908933
transform -1 0 13248 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_7
timestamp 1626908933
transform 1 0 12864 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_6
timestamp 1626908933
transform -1 0 13248 0 1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2621
timestamp 1626908933
transform 1 0 13296 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_686
timestamp 1626908933
transform 1 0 13296 0 1 10545
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2636
timestamp 1626908933
transform 1 0 13200 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_669
timestamp 1626908933
transform 1 0 13200 0 1 10545
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1422
timestamp 1626908933
transform 1 0 13248 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_431
timestamp 1626908933
transform 1 0 13248 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_827
timestamp 1626908933
transform 1 0 13248 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_226
timestamp 1626908933
transform 1 0 13248 0 -1 10656
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1168
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_520
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1168
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_520
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_947
timestamp 1626908933
transform 1 0 13440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_349
timestamp 1626908933
transform 1 0 13440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_444
timestamp 1626908933
transform 1 0 13344 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1166
timestamp 1626908933
transform 1 0 13344 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_33
timestamp 1626908933
transform 1 0 13824 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_8
timestamp 1626908933
transform 1 0 13824 0 -1 10656
box -38 -49 2246 715
use M1M2_PR  M1M2_PR_779
timestamp 1626908933
transform 1 0 14544 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1514
timestamp 1626908933
transform 1 0 13968 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2746
timestamp 1626908933
transform 1 0 14544 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3481
timestamp 1626908933
transform 1 0 13968 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1602
timestamp 1626908933
transform 1 0 13872 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3537
timestamp 1626908933
transform 1 0 13872 0 1 10249
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1667
timestamp 1626908933
transform 1 0 14256 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3634
timestamp 1626908933
transform 1 0 14256 0 1 10397
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1749
timestamp 1626908933
transform 1 0 14160 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3684
timestamp 1626908933
transform 1 0 14160 0 1 10397
box -29 -23 29 23
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_3
timestamp 1626908933
transform -1 0 14688 0 1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_9
timestamp 1626908933
transform -1 0 14688 0 1 10656
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_832
timestamp 1626908933
transform 1 0 14900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_184
timestamp 1626908933
transform 1 0 14900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_832
timestamp 1626908933
transform 1 0 14900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_184
timestamp 1626908933
transform 1 0 14900 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1777
timestamp 1626908933
transform 1 0 14880 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_786
timestamp 1626908933
transform 1 0 14880 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_591
timestamp 1626908933
transform 1 0 14976 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_234
timestamp 1626908933
transform 1 0 14976 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1040
timestamp 1626908933
transform 1 0 14688 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_439
timestamp 1626908933
transform 1 0 14688 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_440
timestamp 1626908933
transform 1 0 15456 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1041
timestamp 1626908933
transform 1 0 15456 0 1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_743
timestamp 1626908933
transform 1 0 15312 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1712
timestamp 1626908933
transform 1 0 15504 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2710
timestamp 1626908933
transform 1 0 15312 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3679
timestamp 1626908933
transform 1 0 15504 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_322
timestamp 1626908933
transform 1 0 15072 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_920
timestamp 1626908933
transform 1 0 15072 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_787
timestamp 1626908933
transform 1 0 15648 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1778
timestamp 1626908933
transform 1 0 15648 0 1 10656
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1144
timestamp 1626908933
transform 1 0 16100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_496
timestamp 1626908933
transform 1 0 16100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1144
timestamp 1626908933
transform 1 0 16100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_496
timestamp 1626908933
transform 1 0 16100 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1421
timestamp 1626908933
transform 1 0 16128 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_430
timestamp 1626908933
transform 1 0 16128 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2560
timestamp 1626908933
transform 1 0 16272 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_593
timestamp 1626908933
transform 1 0 16272 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1767
timestamp 1626908933
transform 1 0 16224 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_776
timestamp 1626908933
transform 1 0 16224 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1034
timestamp 1626908933
transform 1 0 16032 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_433
timestamp 1626908933
transform 1 0 16032 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_101
timestamp 1626908933
transform 1 0 16320 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_32
timestamp 1626908933
transform 1 0 16320 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_393
timestamp 1626908933
transform 1 0 16224 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1115
timestamp 1626908933
transform 1 0 16224 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_9
timestamp 1626908933
transform 1 0 15744 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_71
timestamp 1626908933
transform 1 0 15744 0 1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2700
timestamp 1626908933
transform 1 0 16464 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_765
timestamp 1626908933
transform 1 0 16464 0 1 10545
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_220
timestamp 1626908933
transform 1 0 16992 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_821
timestamp 1626908933
transform 1 0 16992 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_777
timestamp 1626908933
transform 1 0 16800 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1768
timestamp 1626908933
transform 1 0 16800 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_589
timestamp 1626908933
transform 1 0 17040 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_601
timestamp 1626908933
transform 1 0 17040 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2524
timestamp 1626908933
transform 1 0 17040 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2536
timestamp 1626908933
transform 1 0 17040 0 1 10397
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_808
timestamp 1626908933
transform 1 0 17300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_160
timestamp 1626908933
transform 1 0 17300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_808
timestamp 1626908933
transform 1 0 17300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_160
timestamp 1626908933
transform 1 0 17300 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2533
timestamp 1626908933
transform 1 0 17136 0 1 10471
box -29 -23 29 23
use L1M1_PR  L1M1_PR_598
timestamp 1626908933
transform 1 0 17136 0 1 10471
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1420
timestamp 1626908933
transform 1 0 17184 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_429
timestamp 1626908933
transform 1 0 17184 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2532
timestamp 1626908933
transform 1 0 17328 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2530
timestamp 1626908933
transform 1 0 17424 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_597
timestamp 1626908933
transform 1 0 17328 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_595
timestamp 1626908933
transform 1 0 17424 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2555
timestamp 1626908933
transform 1 0 17520 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_588
timestamp 1626908933
transform 1 0 17520 0 1 10101
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_598
timestamp 1626908933
transform 1 0 17472 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_241
timestamp 1626908933
transform 1 0 17472 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_879
timestamp 1626908933
transform 1 0 17280 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_281
timestamp 1626908933
transform 1 0 17280 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_0
timestamp 1626908933
transform -1 0 17472 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_6
timestamp 1626908933
transform -1 0 17472 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_270
timestamp 1626908933
transform 1 0 17664 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_868
timestamp 1626908933
transform 1 0 17664 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_445
timestamp 1626908933
transform 1 0 17568 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1436
timestamp 1626908933
transform 1 0 17568 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_582
timestamp 1626908933
transform 1 0 17712 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_586
timestamp 1626908933
transform 1 0 17808 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2549
timestamp 1626908933
transform 1 0 17712 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2553
timestamp 1626908933
transform 1 0 17808 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_758
timestamp 1626908933
transform 1 0 18192 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2725
timestamp 1626908933
transform 1 0 18192 0 1 10101
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_472
timestamp 1626908933
transform 1 0 18500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1120
timestamp 1626908933
transform 1 0 18500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_472
timestamp 1626908933
transform 1 0 18500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1120
timestamp 1626908933
transform 1 0 18500 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_359
timestamp 1626908933
transform 1 0 18048 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1081
timestamp 1626908933
transform 1 0 18048 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__a31oi_2  sky130_fd_sc_hs__a31oi_2_0
timestamp 1626908933
transform 1 0 17664 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__a31oi_2  sky130_fd_sc_hs__a31oi_2_1
timestamp 1626908933
transform 1 0 17664 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_23
timestamp 1626908933
transform 1 0 18528 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_75
timestamp 1626908933
transform 1 0 18528 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_441
timestamp 1626908933
transform 1 0 18912 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1042
timestamp 1626908933
transform 1 0 18912 0 1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_786
timestamp 1626908933
transform 1 0 18864 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2721
timestamp 1626908933
transform 1 0 18864 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_809
timestamp 1626908933
transform 1 0 19152 0 1 10175
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2744
timestamp 1626908933
transform 1 0 19152 0 1 10175
box -29 -23 29 23
use M1M2_PR  M1M2_PR_681
timestamp 1626908933
transform 1 0 18960 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2648
timestamp 1626908933
transform 1 0 18960 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_693
timestamp 1626908933
transform 1 0 19056 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_698
timestamp 1626908933
transform 1 0 18960 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2628
timestamp 1626908933
transform 1 0 19056 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2633
timestamp 1626908933
transform 1 0 18960 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_788
timestamp 1626908933
transform 1 0 19104 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1779
timestamp 1626908933
transform 1 0 19104 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2464
timestamp 1626908933
transform 1 0 19344 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_529
timestamp 1626908933
transform 1 0 19344 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2642
timestamp 1626908933
transform 1 0 19248 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2495
timestamp 1626908933
transform 1 0 19344 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_675
timestamp 1626908933
transform 1 0 19248 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_528
timestamp 1626908933
transform 1 0 19344 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_70
timestamp 1626908933
transform 1 0 19200 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_8
timestamp 1626908933
transform 1 0 19200 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__nor4_1  sky130_fd_sc_hs__nor4_1_1
timestamp 1626908933
transform -1 0 19392 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__nor4_1  sky130_fd_sc_hs__nor4_1_3
timestamp 1626908933
transform -1 0 19392 0 -1 10656
box -38 -49 614 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_136
timestamp 1626908933
transform 1 0 19700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_784
timestamp 1626908933
transform 1 0 19700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_136
timestamp 1626908933
transform 1 0 19700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_784
timestamp 1626908933
transform 1 0 19700 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_233
timestamp 1626908933
transform 1 0 19968 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_590
timestamp 1626908933
transform 1 0 19968 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_442
timestamp 1626908933
transform 1 0 20064 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1043
timestamp 1626908933
transform 1 0 20064 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_444
timestamp 1626908933
transform 1 0 20160 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1435
timestamp 1626908933
transform 1 0 20160 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_330
timestamp 1626908933
transform 1 0 19392 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1052
timestamp 1626908933
transform 1 0 19392 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_24
timestamp 1626908933
transform 1 0 19584 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_76
timestamp 1626908933
transform 1 0 19584 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_789
timestamp 1626908933
transform 1 0 20256 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1780
timestamp 1626908933
transform 1 0 20256 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_219
timestamp 1626908933
transform 1 0 20736 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_820
timestamp 1626908933
transform 1 0 20736 0 1 10656
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_448
timestamp 1626908933
transform 1 0 20900 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1096
timestamp 1626908933
transform 1 0 20900 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_448
timestamp 1626908933
transform 1 0 20900 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1096
timestamp 1626908933
transform 1 0 20900 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_301
timestamp 1626908933
transform 1 0 20640 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1023
timestamp 1626908933
transform 1 0 20640 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_204
timestamp 1626908933
transform 1 0 20928 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_218
timestamp 1626908933
transform 1 0 20256 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_802
timestamp 1626908933
transform 1 0 20928 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_816
timestamp 1626908933
transform 1 0 20256 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_1
timestamp 1626908933
transform 1 0 20352 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_63
timestamp 1626908933
transform 1 0 20352 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_225
timestamp 1626908933
transform 1 0 21408 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_826
timestamp 1626908933
transform 1 0 21408 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_443
timestamp 1626908933
transform 1 0 21600 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1434
timestamp 1626908933
transform 1 0 21600 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_559
timestamp 1626908933
transform 1 0 21744 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2526
timestamp 1626908933
transform 1 0 21744 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_593
timestamp 1626908933
transform 1 0 21648 0 1 10471
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2528
timestamp 1626908933
transform 1 0 21648 0 1 10471
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_284
timestamp 1626908933
transform 1 0 21312 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1006
timestamp 1626908933
transform 1 0 21312 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_3
timestamp 1626908933
transform 1 0 21696 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  sky130_fd_sc_hs__nor3_1_11
timestamp 1626908933
transform 1 0 21696 0 -1 10656
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_760
timestamp 1626908933
transform 1 0 22100 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_112
timestamp 1626908933
transform 1 0 22100 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_760
timestamp 1626908933
transform 1 0 22100 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_112
timestamp 1626908933
transform 1 0 22100 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2668
timestamp 1626908933
transform 1 0 22032 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_733
timestamp 1626908933
transform 1 0 22032 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2497
timestamp 1626908933
transform 1 0 21936 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_562
timestamp 1626908933
transform 1 0 21936 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_819
timestamp 1626908933
transform 1 0 22080 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_218
timestamp 1626908933
transform 1 0 22080 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_22
timestamp 1626908933
transform 1 0 22080 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_74
timestamp 1626908933
transform 1 0 22080 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_240
timestamp 1626908933
transform 1 0 22464 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_597
timestamp 1626908933
transform 1 0 22464 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_710
timestamp 1626908933
transform 1 0 22320 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2677
timestamp 1626908933
transform 1 0 22320 0 1 10101
box -32 -32 32 32
use L1M1_PR  L1M1_PR_559
timestamp 1626908933
transform 1 0 22128 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2494
timestamp 1626908933
transform 1 0 22128 0 1 10249
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_251
timestamp 1626908933
transform 1 0 22272 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_252
timestamp 1626908933
transform 1 0 22560 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_973
timestamp 1626908933
transform 1 0 22272 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_974
timestamp 1626908933
transform 1 0 22560 0 -1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2534
timestamp 1626908933
transform 1 0 23280 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_567
timestamp 1626908933
transform 1 0 23280 0 1 10101
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1072
timestamp 1626908933
transform 1 0 23300 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_424
timestamp 1626908933
transform 1 0 23300 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1072
timestamp 1626908933
transform 1 0 23300 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_424
timestamp 1626908933
transform 1 0 23300 0 1 10656
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2529
timestamp 1626908933
transform 1 0 23088 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_562
timestamp 1626908933
transform 1 0 23088 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1035
timestamp 1626908933
transform 1 0 23328 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_434
timestamp 1626908933
transform 1 0 23328 0 -1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_2528
timestamp 1626908933
transform 1 0 23472 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_561
timestamp 1626908933
transform 1 0 23472 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1769
timestamp 1626908933
transform 1 0 23520 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_778
timestamp 1626908933
transform 1 0 23520 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2505
timestamp 1626908933
transform 1 0 23568 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_570
timestamp 1626908933
transform 1 0 23568 0 1 10101
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2517
timestamp 1626908933
transform 1 0 23664 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_550
timestamp 1626908933
transform 1 0 23664 0 1 10101
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2499
timestamp 1626908933
transform 1 0 23760 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_564
timestamp 1626908933
transform 1 0 23760 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2533
timestamp 1626908933
transform 1 0 23760 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_566
timestamp 1626908933
transform 1 0 23760 0 1 10175
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_93
timestamp 1626908933
transform -1 0 23520 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_24
timestamp 1626908933
transform -1 0 23520 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_12
timestamp 1626908933
transform 1 0 23520 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_35
timestamp 1626908933
transform 1 0 23520 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_0
timestamp 1626908933
transform -1 0 24192 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_4
timestamp 1626908933
transform -1 0 24192 0 -1 10656
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2490
timestamp 1626908933
transform 1 0 23856 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_555
timestamp 1626908933
transform 1 0 23856 0 1 10101
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2519
timestamp 1626908933
transform 1 0 23856 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_552
timestamp 1626908933
transform 1 0 23856 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2496
timestamp 1626908933
transform 1 0 24048 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2027
timestamp 1626908933
transform 1 0 24144 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_561
timestamp 1626908933
transform 1 0 24048 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_92
timestamp 1626908933
transform 1 0 24144 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2522
timestamp 1626908933
transform 1 0 24048 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_555
timestamp 1626908933
transform 1 0 24048 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_825
timestamp 1626908933
transform 1 0 24192 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_224
timestamp 1626908933
transform 1 0 24192 0 -1 10656
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_736
timestamp 1626908933
transform 1 0 24500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_88
timestamp 1626908933
transform 1 0 24500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_736
timestamp 1626908933
transform 1 0 24500 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_88
timestamp 1626908933
transform 1 0 24500 0 1 9990
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2050
timestamp 1626908933
transform 1 0 24240 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_83
timestamp 1626908933
transform 1 0 24240 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1433
timestamp 1626908933
transform 1 0 24384 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_442
timestamp 1626908933
transform 1 0 24384 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_69
timestamp 1626908933
transform -1 0 24576 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_7
timestamp 1626908933
transform -1 0 24576 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_204
timestamp 1626908933
transform 1 0 24480 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_926
timestamp 1626908933
transform 1 0 24480 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_25
timestamp 1626908933
transform 1 0 24576 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_77
timestamp 1626908933
transform 1 0 24576 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_232
timestamp 1626908933
transform 1 0 24960 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_589
timestamp 1626908933
transform 1 0 24960 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_117
timestamp 1626908933
transform 1 0 25440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_715
timestamp 1626908933
transform 1 0 25440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_223
timestamp 1626908933
transform 1 0 25248 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_824
timestamp 1626908933
transform 1 0 25248 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_428
timestamp 1626908933
transform 1 0 25056 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1419
timestamp 1626908933
transform 1 0 25056 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_754
timestamp 1626908933
transform 1 0 25872 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2689
timestamp 1626908933
transform 1 0 25872 0 1 10545
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_400
timestamp 1626908933
transform 1 0 25700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1048
timestamp 1626908933
transform 1 0 25700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_400
timestamp 1626908933
transform 1 0 25700 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1048
timestamp 1626908933
transform 1 0 25700 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_427
timestamp 1626908933
transform 1 0 25920 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_441
timestamp 1626908933
transform 1 0 25824 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1418
timestamp 1626908933
transform 1 0 25920 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1432
timestamp 1626908933
transform 1 0 25824 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_790
timestamp 1626908933
transform 1 0 26016 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1781
timestamp 1626908933
transform 1 0 26016 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_730
timestamp 1626908933
transform 1 0 26064 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2697
timestamp 1626908933
transform 1 0 26064 0 1 10545
box -32 -32 32 32
use L1M1_PR  L1M1_PR_557
timestamp 1626908933
transform 1 0 25968 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2492
timestamp 1626908933
transform 1 0 25968 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_102
timestamp 1626908933
transform 1 0 26256 0 1 10471
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2037
timestamp 1626908933
transform 1 0 26256 0 1 10471
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_222
timestamp 1626908933
transform 1 0 26208 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_823
timestamp 1626908933
transform 1 0 26208 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_68
timestamp 1626908933
transform -1 0 26208 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_6
timestamp 1626908933
transform -1 0 26208 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_70
timestamp 1626908933
transform 1 0 26112 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_9
timestamp 1626908933
transform 1 0 26112 0 1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_190
timestamp 1626908933
transform 1 0 25152 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_912
timestamp 1626908933
transform 1 0 25152 0 1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2058
timestamp 1626908933
transform 1 0 26448 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_91
timestamp 1626908933
transform 1 0 26448 0 1 10471
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1431
timestamp 1626908933
transform 1 0 26400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1417
timestamp 1626908933
transform 1 0 26400 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_440
timestamp 1626908933
transform 1 0 26400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_426
timestamp 1626908933
transform 1 0 26400 0 1 10656
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_712
timestamp 1626908933
transform 1 0 26900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_64
timestamp 1626908933
transform 1 0 26900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_712
timestamp 1626908933
transform 1 0 26900 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_64
timestamp 1626908933
transform 1 0 26900 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1430
timestamp 1626908933
transform 1 0 27264 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1416
timestamp 1626908933
transform 1 0 27264 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_439
timestamp 1626908933
transform 1 0 27264 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_425
timestamp 1626908933
transform 1 0 27264 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3467
timestamp 1626908933
transform 1 0 27600 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1532
timestamp 1626908933
transform 1 0 27600 0 1 10249
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3619
timestamp 1626908933
transform 1 0 27408 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1652
timestamp 1626908933
transform 1 0 27408 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1770
timestamp 1626908933
transform 1 0 27360 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_779
timestamp 1626908933
transform 1 0 27360 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_596
timestamp 1626908933
transform 1 0 27456 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_239
timestamp 1626908933
transform 1 0 27456 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_684
timestamp 1626908933
transform 1 0 27360 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_86
timestamp 1626908933
transform 1 0 27360 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_161
timestamp 1626908933
transform 1 0 26496 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_162
timestamp 1626908933
transform 1 0 26496 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_883
timestamp 1626908933
transform 1 0 26496 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_884
timestamp 1626908933
transform 1 0 26496 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_41
timestamp 1626908933
transform 1 0 27552 0 -1 10656
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_17
timestamp 1626908933
transform 1 0 27552 0 -1 10656
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_1446
timestamp 1626908933
transform 1 0 27696 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1678
timestamp 1626908933
transform 1 0 27888 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3413
timestamp 1626908933
transform 1 0 27696 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3645
timestamp 1626908933
transform 1 0 27888 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1733
timestamp 1626908933
transform 1 0 27984 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3668
timestamp 1626908933
transform 1 0 27984 0 1 10323
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_376
timestamp 1626908933
transform 1 0 28100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1024
timestamp 1626908933
transform 1 0 28100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_376
timestamp 1626908933
transform 1 0 28100 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1024
timestamp 1626908933
transform 1 0 28100 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_128
timestamp 1626908933
transform 1 0 27744 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_850
timestamp 1626908933
transform 1 0 27744 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_424
timestamp 1626908933
transform 1 0 28896 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1415
timestamp 1626908933
transform 1 0 28896 0 1 10656
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_40
timestamp 1626908933
transform 1 0 29300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_688
timestamp 1626908933
transform 1 0 29300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_40
timestamp 1626908933
transform 1 0 29300 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_688
timestamp 1626908933
transform 1 0 29300 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_93
timestamp 1626908933
transform 1 0 28992 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_815
timestamp 1626908933
transform 1 0 28992 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_63
timestamp 1626908933
transform 1 0 28512 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_661
timestamp 1626908933
transform 1 0 28512 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_423
timestamp 1626908933
transform 1 0 29760 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1414
timestamp 1626908933
transform 1 0 29760 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_88
timestamp 1626908933
transform 1 0 29520 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2055
timestamp 1626908933
transform 1 0 29520 0 1 10471
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2034
timestamp 1626908933
transform 1 0 29808 0 1 10471
box -29 -23 29 23
use L1M1_PR  L1M1_PR_99
timestamp 1626908933
transform 1 0 29808 0 1 10471
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1782
timestamp 1626908933
transform 1 0 29856 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1429
timestamp 1626908933
transform 1 0 29856 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_791
timestamp 1626908933
transform 1 0 29856 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_438
timestamp 1626908933
transform 1 0 29856 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_588
timestamp 1626908933
transform 1 0 29952 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_231
timestamp 1626908933
transform 1 0 29952 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_818
timestamp 1626908933
transform 1 0 30048 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_217
timestamp 1626908933
transform 1 0 30048 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_31
timestamp 1626908933
transform 1 0 29952 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_629
timestamp 1626908933
transform 1 0 29952 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1413
timestamp 1626908933
transform 1 0 30240 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_422
timestamp 1626908933
transform 1 0 30240 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_775
timestamp 1626908933
transform 1 0 30336 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_774
timestamp 1626908933
transform 1 0 30336 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_53
timestamp 1626908933
transform 1 0 30336 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_52
timestamp 1626908933
transform 1 0 30336 0 1 10656
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_352
timestamp 1626908933
transform 1 0 30500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1000
timestamp 1626908933
transform 1 0 30500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_352
timestamp 1626908933
transform 1 0 30500 0 1 10656
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1000
timestamp 1626908933
transform 1 0 30500 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_421
timestamp 1626908933
transform 1 0 31104 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1412
timestamp 1626908933
transform 1 0 31104 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_15
timestamp 1626908933
transform 1 0 31200 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_737
timestamp 1626908933
transform 1 0 31200 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_9
timestamp 1626908933
transform 1 0 31104 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_607
timestamp 1626908933
transform 1 0 31104 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_437
timestamp 1626908933
transform 1 0 31488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1428
timestamp 1626908933
transform 1 0 31488 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1792
timestamp 1626908933
transform 1 0 31344 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3759
timestamp 1626908933
transform 1 0 31344 0 1 10471
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_664
timestamp 1626908933
transform 1 0 31700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_16
timestamp 1626908933
transform 1 0 31700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_664
timestamp 1626908933
transform 1 0 31700 0 1 9990
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_16
timestamp 1626908933
transform 1 0 31700 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1771
timestamp 1626908933
transform 1 0 31584 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_780
timestamp 1626908933
transform 1 0 31584 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1036
timestamp 1626908933
transform 1 0 31776 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_435
timestamp 1626908933
transform 1 0 31776 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_595
timestamp 1626908933
transform 1 0 31680 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_238
timestamp 1626908933
transform 1 0 31680 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_781
timestamp 1626908933
transform 1 0 31968 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_792
timestamp 1626908933
transform 1 0 31968 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1772
timestamp 1626908933
transform 1 0 31968 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1783
timestamp 1626908933
transform 1 0 31968 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1790
timestamp 1626908933
transform 1 0 32016 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3757
timestamp 1626908933
transform 1 0 32016 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3870
timestamp 1626908933
transform 1 0 48 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1903
timestamp 1626908933
transform 1 0 48 0 1 10989
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1411
timestamp 1626908933
transform 1 0 0 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_420
timestamp 1626908933
transform 1 0 0 0 -1 11988
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_975
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_327
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_975
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_327
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1194
timestamp 1626908933
transform 1 0 96 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_596
timestamp 1626908933
transform 1 0 96 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_419
timestamp 1626908933
transform 1 0 1344 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1410
timestamp 1626908933
transform 1 0 1344 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1767
timestamp 1626908933
transform 1 0 1104 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3734
timestamp 1626908933
transform 1 0 1104 0 1 10767
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1398
timestamp 1626908933
transform 1 0 1296 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1783
timestamp 1626908933
transform 1 0 1008 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3333
timestamp 1626908933
transform 1 0 1296 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3718
timestamp 1626908933
transform 1 0 1008 0 1 10767
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_4
timestamp 1626908933
transform 1 0 480 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_12
timestamp 1626908933
transform 1 0 480 0 -1 11988
box -38 -49 902 715
use M1M2_PR  M1M2_PR_312
timestamp 1626908933
transform 1 0 1968 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1318
timestamp 1626908933
transform 1 0 1392 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2279
timestamp 1626908933
transform 1 0 1968 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3285
timestamp 1626908933
transform 1 0 1392 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1414
timestamp 1626908933
transform 1 0 1392 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3349
timestamp 1626908933
transform 1 0 1392 0 1 10767
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_817
timestamp 1626908933
transform 1 0 2208 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_216
timestamp 1626908933
transform 1 0 2208 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3301
timestamp 1626908933
transform 1 0 2448 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1334
timestamp 1626908933
transform 1 0 2448 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1409
timestamp 1626908933
transform 1 0 2400 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_418
timestamp 1626908933
transform 1 0 2400 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_587
timestamp 1626908933
transform 1 0 2496 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_230
timestamp 1626908933
transform 1 0 2496 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2274
timestamp 1626908933
transform 1 0 2736 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_339
timestamp 1626908933
transform 1 0 2736 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_681
timestamp 1626908933
transform 1 0 1440 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1403
timestamp 1626908933
transform 1 0 1440 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_8
timestamp 1626908933
transform -1 0 4320 0 -1 11988
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_2
timestamp 1626908933
transform -1 0 4320 0 -1 11988
box -38 -49 1766 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_951
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_303
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_951
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_303
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2293
timestamp 1626908933
transform 1 0 3216 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_358
timestamp 1626908933
transform 1 0 3216 0 1 10767
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2297
timestamp 1626908933
transform 1 0 3696 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_330
timestamp 1626908933
transform 1 0 3696 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_520
timestamp 1626908933
transform 1 0 4512 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1118
timestamp 1626908933
transform 1 0 4512 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_215
timestamp 1626908933
transform 1 0 4320 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_816
timestamp 1626908933
transform 1 0 4320 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1325
timestamp 1626908933
transform 1 0 4368 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3292
timestamp 1626908933
transform 1 0 4368 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1406
timestamp 1626908933
transform 1 0 4368 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3341
timestamp 1626908933
transform 1 0 4368 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_317
timestamp 1626908933
transform 1 0 4656 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1390
timestamp 1626908933
transform 1 0 4848 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2284
timestamp 1626908933
transform 1 0 4656 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3357
timestamp 1626908933
transform 1 0 4848 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_343
timestamp 1626908933
transform 1 0 5040 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1471
timestamp 1626908933
transform 1 0 4848 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2278
timestamp 1626908933
transform 1 0 5040 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3406
timestamp 1626908933
transform 1 0 4848 0 1 11211
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_279
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_927
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_279
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_927
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_10
timestamp 1626908933
transform -1 0 6624 0 -1 11988
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_4
timestamp 1626908933
transform -1 0 6624 0 -1 11988
box -38 -49 1766 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_87
timestamp 1626908933
transform -1 0 7392 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_25
timestamp 1626908933
transform -1 0 7392 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1079
timestamp 1626908933
transform 1 0 6624 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_481
timestamp 1626908933
transform 1 0 6624 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1784
timestamp 1626908933
transform 1 0 7392 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_793
timestamp 1626908933
transform 1 0 7392 0 -1 11988
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_903
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_255
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_903
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_255
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_586
timestamp 1626908933
transform 1 0 7488 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_229
timestamp 1626908933
transform 1 0 7488 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_815
timestamp 1626908933
transform 1 0 7584 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_214
timestamp 1626908933
transform 1 0 7584 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_417
timestamp 1626908933
transform 1 0 7776 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1408
timestamp 1626908933
transform 1 0 7776 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_840
timestamp 1626908933
transform 1 0 8016 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2775
timestamp 1626908933
transform 1 0 8016 0 1 11211
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_557
timestamp 1626908933
transform 1 0 7872 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1279
timestamp 1626908933
transform 1 0 7872 0 -1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2779
timestamp 1626908933
transform 1 0 8208 0 1 11137
box -29 -23 29 23
use L1M1_PR  L1M1_PR_844
timestamp 1626908933
transform 1 0 8208 0 1 11137
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2773
timestamp 1626908933
transform 1 0 8112 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_806
timestamp 1626908933
transform 1 0 8112 0 1 11211
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_416
timestamp 1626908933
transform 1 0 8640 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1407
timestamp 1626908933
transform 1 0 8640 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1480
timestamp 1626908933
transform 1 0 8688 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3447
timestamp 1626908933
transform 1 0 8688 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_803
timestamp 1626908933
transform 1 0 8880 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_809
timestamp 1626908933
transform 1 0 9072 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2770
timestamp 1626908933
transform 1 0 8880 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2776
timestamp 1626908933
transform 1 0 9072 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_837
timestamp 1626908933
transform 1 0 8880 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1567
timestamp 1626908933
transform 1 0 9072 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2772
timestamp 1626908933
transform 1 0 8880 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3502
timestamp 1626908933
transform 1 0 9072 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_538
timestamp 1626908933
transform 1 0 9120 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1260
timestamp 1626908933
transform 1 0 9120 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_13
timestamp 1626908933
transform 1 0 8736 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_75
timestamp 1626908933
transform 1 0 8736 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1955
timestamp 1626908933
transform 1 0 9936 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_20
timestamp 1626908933
transform 1 0 9936 0 1 10767
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1986
timestamp 1626908933
transform 1 0 9936 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_19
timestamp 1626908933
transform 1 0 9936 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1406
timestamp 1626908933
transform 1 0 9888 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_415
timestamp 1626908933
transform 1 0 9888 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1021
timestamp 1626908933
transform 1 0 9984 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_423
timestamp 1626908933
transform 1 0 9984 0 -1 11988
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_879
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_231
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_879
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_231
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_55
timestamp 1626908933
transform 1 0 10368 0 -1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_16
timestamp 1626908933
transform 1 0 10368 0 -1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1405
timestamp 1626908933
transform 1 0 10944 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_414
timestamp 1626908933
transform 1 0 10944 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1218
timestamp 1626908933
transform 1 0 11040 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_496
timestamp 1626908933
transform 1 0 11040 0 -1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_666
timestamp 1626908933
transform 1 0 11472 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2633
timestamp 1626908933
transform 1 0 11472 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_213
timestamp 1626908933
transform 1 0 11808 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_814
timestamp 1626908933
transform 1 0 11808 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_63
timestamp 1626908933
transform 1 0 11760 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2030
timestamp 1626908933
transform 1 0 11760 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_70
timestamp 1626908933
transform 1 0 11856 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_683
timestamp 1626908933
transform 1 0 11760 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2005
timestamp 1626908933
transform 1 0 11856 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2618
timestamp 1626908933
transform 1 0 11760 0 1 10767
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_413
timestamp 1626908933
transform 1 0 12000 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1404
timestamp 1626908933
transform 1 0 12000 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_153
timestamp 1626908933
transform 1 0 12048 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2120
timestamp 1626908933
transform 1 0 12048 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_169
timestamp 1626908933
transform 1 0 12048 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2104
timestamp 1626908933
transform 1 0 12048 0 1 10915
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_228
timestamp 1626908933
transform 1 0 12480 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_585
timestamp 1626908933
transform 1 0 12480 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_682
timestamp 1626908933
transform 1 0 12720 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2617
timestamp 1626908933
transform 1 0 12720 0 1 10767
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_207
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_855
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_207
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_855
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_462
timestamp 1626908933
transform 1 0 12576 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1184
timestamp 1626908933
transform 1 0 12576 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_379
timestamp 1626908933
transform 1 0 12096 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_977
timestamp 1626908933
transform 1 0 12096 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_590
timestamp 1626908933
transform 1 0 13008 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_664
timestamp 1626908933
transform 1 0 13392 0 1 10841
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2557
timestamp 1626908933
transform 1 0 13008 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2631
timestamp 1626908933
transform 1 0 13392 0 1 10841
box -32 -32 32 32
use L1M1_PR  L1M1_PR_599
timestamp 1626908933
transform 1 0 13104 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_681
timestamp 1626908933
transform 1 0 13296 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2534
timestamp 1626908933
transform 1 0 13104 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2616
timestamp 1626908933
transform 1 0 13296 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_663
timestamp 1626908933
transform 1 0 12912 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_668
timestamp 1626908933
transform 1 0 13200 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2630
timestamp 1626908933
transform 1 0 12912 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2635
timestamp 1626908933
transform 1 0 13200 0 1 11433
box -32 -32 32 32
use L1M1_PR  L1M1_PR_678
timestamp 1626908933
transform 1 0 12912 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_685
timestamp 1626908933
transform 1 0 13584 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2613
timestamp 1626908933
transform 1 0 12912 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2620
timestamp 1626908933
transform 1 0 13584 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__o2bb2ai_1  sky130_fd_sc_hs__o2bb2ai_1_0
timestamp 1626908933
transform -1 0 14016 0 -1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__o2bb2ai_1  sky130_fd_sc_hs__o2bb2ai_1_1
timestamp 1626908933
transform -1 0 14016 0 -1 11988
box -38 -49 710 715
use M1M2_PR  M1M2_PR_2736
timestamp 1626908933
transform 1 0 13776 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_769
timestamp 1626908933
transform 1 0 13776 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1995
timestamp 1626908933
transform 1 0 14064 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_60
timestamp 1626908933
transform 1 0 14064 0 1 11211
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2022
timestamp 1626908933
transform 1 0 14064 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_55
timestamp 1626908933
transform 1 0 14064 0 1 11211
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1403
timestamp 1626908933
transform 1 0 14016 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_412
timestamp 1626908933
transform 1 0 14016 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2734
timestamp 1626908933
transform 1 0 14352 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2703
timestamp 1626908933
transform 1 0 14448 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_799
timestamp 1626908933
transform 1 0 14352 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_768
timestamp 1626908933
transform 1 0 14448 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2614
timestamp 1626908933
transform 1 0 14544 0 1 10841
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1991
timestamp 1626908933
transform 1 0 14640 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_679
timestamp 1626908933
transform 1 0 14544 0 1 10841
box -29 -23 29 23
use L1M1_PR  L1M1_PR_56
timestamp 1626908933
transform 1 0 14640 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2017
timestamp 1626908933
transform 1 0 14736 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_50
timestamp 1626908933
transform 1 0 14736 0 1 10915
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_831
timestamp 1626908933
transform 1 0 14900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_183
timestamp 1626908933
transform 1 0 14900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_831
timestamp 1626908933
transform 1 0 14900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_183
timestamp 1626908933
transform 1 0 14900 0 1 11322
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2016
timestamp 1626908933
transform 1 0 14736 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_49
timestamp 1626908933
transform 1 0 14736 0 1 11433
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1990
timestamp 1626908933
transform 1 0 14928 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_55
timestamp 1626908933
transform 1 0 14928 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_431
timestamp 1626908933
transform 1 0 14112 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1153
timestamp 1626908933
transform 1 0 14112 0 -1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_603
timestamp 1626908933
transform 1 0 15984 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2538
timestamp 1626908933
transform 1 0 15984 0 1 10767
box -29 -23 29 23
use M1M2_PR  M1M2_PR_592
timestamp 1626908933
transform 1 0 16272 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_746
timestamp 1626908933
transform 1 0 16272 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2559
timestamp 1626908933
transform 1 0 16272 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2713
timestamp 1626908933
transform 1 0 16272 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_771
timestamp 1626908933
transform 1 0 16080 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2706
timestamp 1626908933
transform 1 0 16080 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_742
timestamp 1626908933
transform 1 0 15312 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2709
timestamp 1626908933
transform 1 0 15312 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_766
timestamp 1626908933
transform 1 0 15696 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2701
timestamp 1626908933
transform 1 0 15696 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_53
timestamp 1626908933
transform 1 0 15888 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1988
timestamp 1626908933
transform 1 0 15888 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_32
timestamp 1626908933
transform -1 0 17184 0 -1 11988
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_8
timestamp 1626908933
transform -1 0 17184 0 -1 11988
box -38 -49 2342 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_807
timestamp 1626908933
transform 1 0 17300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_159
timestamp 1626908933
transform 1 0 17300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_807
timestamp 1626908933
transform 1 0 17300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_159
timestamp 1626908933
transform 1 0 17300 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1785
timestamp 1626908933
transform 1 0 17376 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_794
timestamp 1626908933
transform 1 0 17376 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1044
timestamp 1626908933
transform 1 0 17184 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_443
timestamp 1626908933
transform 1 0 17184 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1402
timestamp 1626908933
transform 1 0 17568 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_411
timestamp 1626908933
transform 1 0 17568 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_584
timestamp 1626908933
transform 1 0 17472 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_227
timestamp 1626908933
transform 1 0 17472 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2523
timestamp 1626908933
transform 1 0 17712 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_588
timestamp 1626908933
transform 1 0 17712 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3869
timestamp 1626908933
transform 1 0 17712 0 1 11137
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2548
timestamp 1626908933
transform 1 0 17712 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1902
timestamp 1626908933
transform 1 0 17712 0 1 11137
box -32 -32 32 32
use M1M2_PR  M1M2_PR_581
timestamp 1626908933
transform 1 0 17712 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2522
timestamp 1626908933
transform 1 0 17808 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_587
timestamp 1626908933
transform 1 0 17808 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_410
timestamp 1626908933
transform 1 0 18048 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1401
timestamp 1626908933
transform 1 0 18048 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_585
timestamp 1626908933
transform 1 0 18096 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2552
timestamp 1626908933
transform 1 0 18096 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_591
timestamp 1626908933
transform 1 0 18192 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2526
timestamp 1626908933
transform 1 0 18192 0 1 10915
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_358
timestamp 1626908933
transform 1 0 18144 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1080
timestamp 1626908933
transform 1 0 18144 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_269
timestamp 1626908933
transform 1 0 17664 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_867
timestamp 1626908933
transform 1 0 17664 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_580
timestamp 1626908933
transform 1 0 18288 0 1 11063
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2547
timestamp 1626908933
transform 1 0 18288 0 1 11063
box -32 -32 32 32
use L1M1_PR  L1M1_PR_531
timestamp 1626908933
transform 1 0 18480 0 1 10841
box -29 -23 29 23
use L1M1_PR  L1M1_PR_585
timestamp 1626908933
transform 1 0 18672 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2466
timestamp 1626908933
transform 1 0 18480 0 1 10841
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2520
timestamp 1626908933
transform 1 0 18672 0 1 11211
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_409
timestamp 1626908933
transform 1 0 18912 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1400
timestamp 1626908933
transform 1 0 18912 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_680
timestamp 1626908933
transform 1 0 18960 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2647
timestamp 1626908933
transform 1 0 18960 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_241
timestamp 1626908933
transform 1 0 19008 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_839
timestamp 1626908933
transform 1 0 19008 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2629
timestamp 1626908933
transform 1 0 19152 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2626
timestamp 1626908933
transform 1 0 19344 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_694
timestamp 1626908933
transform 1 0 19152 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_691
timestamp 1626908933
transform 1 0 19344 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2643
timestamp 1626908933
transform 1 0 19152 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2641
timestamp 1626908933
transform 1 0 19248 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_676
timestamp 1626908933
transform 1 0 19152 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_674
timestamp 1626908933
transform 1 0 19248 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_584
timestamp 1626908933
transform 1 0 19536 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_696
timestamp 1626908933
transform 1 0 19632 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2519
timestamp 1626908933
transform 1 0 19536 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2631
timestamp 1626908933
transform 1 0 19632 0 1 10767
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_135
timestamp 1626908933
transform 1 0 19700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_783
timestamp 1626908933
transform 1 0 19700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_135
timestamp 1626908933
transform 1 0 19700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_783
timestamp 1626908933
transform 1 0 19700 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_408
timestamp 1626908933
transform 1 0 20160 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1399
timestamp 1626908933
transform 1 0 20160 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_679
timestamp 1626908933
transform 1 0 19920 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2646
timestamp 1626908933
transform 1 0 19920 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_329
timestamp 1626908933
transform 1 0 19392 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1051
timestamp 1626908933
transform 1 0 19392 0 -1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2491
timestamp 1626908933
transform 1 0 20496 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_524
timestamp 1626908933
transform 1 0 20496 0 1 10767
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2457
timestamp 1626908933
transform 1 0 20592 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_522
timestamp 1626908933
transform 1 0 20592 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2465
timestamp 1626908933
transform 1 0 20496 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_530
timestamp 1626908933
transform 1 0 20496 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2468
timestamp 1626908933
transform 1 0 20304 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_533
timestamp 1626908933
transform 1 0 20304 0 1 11211
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2498
timestamp 1626908933
transform 1 0 20400 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_531
timestamp 1626908933
transform 1 0 20400 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2467
timestamp 1626908933
transform 1 0 20400 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_532
timestamp 1626908933
transform 1 0 20400 0 1 11433
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2497
timestamp 1626908933
transform 1 0 20400 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_530
timestamp 1626908933
transform 1 0 20400 0 1 11433
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2498
timestamp 1626908933
transform 1 0 20784 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2470
timestamp 1626908933
transform 1 0 20688 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_563
timestamp 1626908933
transform 1 0 20784 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_535
timestamp 1626908933
transform 1 0 20688 0 1 10915
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1786
timestamp 1626908933
transform 1 0 20928 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_795
timestamp 1626908933
transform 1 0 20928 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1045
timestamp 1626908933
transform 1 0 20736 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_444
timestamp 1626908933
transform 1 0 20736 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_76
timestamp 1626908933
transform -1 0 21312 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_15
timestamp 1626908933
transform -1 0 21312 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_72
timestamp 1626908933
transform -1 0 20736 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_3
timestamp 1626908933
transform -1 0 20736 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_407
timestamp 1626908933
transform 1 0 21312 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1398
timestamp 1626908933
transform 1 0 21312 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_532
timestamp 1626908933
transform 1 0 21072 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2499
timestamp 1626908933
transform 1 0 21072 0 1 10915
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_406
timestamp 1626908933
transform 1 0 21792 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1397
timestamp 1626908933
transform 1 0 21792 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_558
timestamp 1626908933
transform 1 0 21744 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2525
timestamp 1626908933
transform 1 0 21744 0 1 11433
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_197
timestamp 1626908933
transform 1 0 21408 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_795
timestamp 1626908933
transform 1 0 21408 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_3
timestamp 1626908933
transform -1 0 22464 0 -1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__o211ai_1  sky130_fd_sc_hs__o211ai_1_9
timestamp 1626908933
transform -1 0 22464 0 -1 11988
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_759
timestamp 1626908933
transform 1 0 22100 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_111
timestamp 1626908933
transform 1 0 22100 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_759
timestamp 1626908933
transform 1 0 22100 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_111
timestamp 1626908933
transform 1 0 22100 0 1 11322
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2753
timestamp 1626908933
transform 1 0 22416 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2515
timestamp 1626908933
transform 1 0 22512 0 1 11063
box -32 -32 32 32
use M1M2_PR  M1M2_PR_786
timestamp 1626908933
transform 1 0 22416 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_548
timestamp 1626908933
transform 1 0 22512 0 1 11063
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_972
timestamp 1626908933
transform 1 0 22560 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_250
timestamp 1626908933
transform 1 0 22560 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_583
timestamp 1626908933
transform 1 0 22464 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_226
timestamp 1626908933
transform 1 0 22464 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_212
timestamp 1626908933
transform 1 0 23328 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_813
timestamp 1626908933
transform 1 0 23328 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_556
timestamp 1626908933
transform 1 0 23280 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_557
timestamp 1626908933
transform 1 0 23280 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2523
timestamp 1626908933
transform 1 0 23280 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2524
timestamp 1626908933
transform 1 0 23280 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_817
timestamp 1626908933
transform 1 0 23184 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2752
timestamp 1626908933
transform 1 0 23184 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_93
timestamp 1626908933
transform 1 0 23568 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2028
timestamp 1626908933
transform 1 0 23568 0 1 10767
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_160
timestamp 1626908933
transform 1 0 23520 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_758
timestamp 1626908933
transform 1 0 23520 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_82
timestamp 1626908933
transform 1 0 24240 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_174
timestamp 1626908933
transform 1 0 24336 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2049
timestamp 1626908933
transform 1 0 24240 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2141
timestamp 1626908933
transform 1 0 24336 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_188
timestamp 1626908933
transform 1 0 24336 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2123
timestamp 1626908933
transform 1 0 24336 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2521
timestamp 1626908933
transform 1 0 24048 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_554
timestamp 1626908933
transform 1 0 24048 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2495
timestamp 1626908933
transform 1 0 24336 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_560
timestamp 1626908933
transform 1 0 24336 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2672
timestamp 1626908933
transform 1 0 24624 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_737
timestamp 1626908933
transform 1 0 24624 0 1 11211
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_735
timestamp 1626908933
transform 1 0 24500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_87
timestamp 1626908933
transform 1 0 24500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_735
timestamp 1626908933
transform 1 0 24500 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_87
timestamp 1626908933
transform 1 0 24500 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_221
timestamp 1626908933
transform 1 0 23904 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_943
timestamp 1626908933
transform 1 0 23904 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1396
timestamp 1626908933
transform 1 0 24672 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_405
timestamp 1626908933
transform 1 0 24672 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_733
timestamp 1626908933
transform 1 0 24768 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_135
timestamp 1626908933
transform 1 0 24768 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2682
timestamp 1626908933
transform 1 0 25008 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_715
timestamp 1626908933
transform 1 0 25008 0 1 11211
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_911
timestamp 1626908933
transform 1 0 25152 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_189
timestamp 1626908933
transform 1 0 25152 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_211
timestamp 1626908933
transform 1 0 25920 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_812
timestamp 1626908933
transform 1 0 25920 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_729
timestamp 1626908933
transform 1 0 26064 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2696
timestamp 1626908933
transform 1 0 26064 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_90
timestamp 1626908933
transform 1 0 26448 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2057
timestamp 1626908933
transform 1 0 26448 0 1 10767
box -32 -32 32 32
use L1M1_PR  L1M1_PR_101
timestamp 1626908933
transform 1 0 26448 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_552
timestamp 1626908933
transform 1 0 26256 0 1 11063
box -29 -23 29 23
use L1M1_PR  L1M1_PR_752
timestamp 1626908933
transform 1 0 26160 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2036
timestamp 1626908933
transform 1 0 26448 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2487
timestamp 1626908933
transform 1 0 26256 0 1 11063
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2687
timestamp 1626908933
transform 1 0 26160 0 1 10915
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_160
timestamp 1626908933
transform 1 0 26496 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_882
timestamp 1626908933
transform 1 0 26496 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_107
timestamp 1626908933
transform 1 0 26112 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_705
timestamp 1626908933
transform 1 0 26112 0 -1 11988
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_711
timestamp 1626908933
transform 1 0 26900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_63
timestamp 1626908933
transform 1 0 26900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_711
timestamp 1626908933
transform 1 0 26900 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_63
timestamp 1626908933
transform 1 0 26900 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1787
timestamp 1626908933
transform 1 0 27360 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1395
timestamp 1626908933
transform 1 0 27264 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_796
timestamp 1626908933
transform 1 0 27360 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_404
timestamp 1626908933
transform 1 0 27264 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_78
timestamp 1626908933
transform 1 0 27552 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_26
timestamp 1626908933
transform 1 0 27552 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_582
timestamp 1626908933
transform 1 0 27456 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_225
timestamp 1626908933
transform 1 0 27456 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_14
timestamp 1626908933
transform 1 0 27936 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_75
timestamp 1626908933
transform 1 0 27936 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_210
timestamp 1626908933
transform 1 0 28224 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_811
timestamp 1626908933
transform 1 0 28224 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_872
timestamp 1626908933
transform 1 0 28272 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2839
timestamp 1626908933
transform 1 0 28272 0 1 11433
box -32 -32 32 32
use L1M1_PR  L1M1_PR_920
timestamp 1626908933
transform 1 0 28080 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2855
timestamp 1626908933
transform 1 0 28080 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_108
timestamp 1626908933
transform 1 0 28416 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_830
timestamp 1626908933
transform 1 0 28416 0 -1 11988
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_687
timestamp 1626908933
transform 1 0 29300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_39
timestamp 1626908933
transform 1 0 29300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_687
timestamp 1626908933
transform 1 0 29300 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_39
timestamp 1626908933
transform 1 0 29300 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_645
timestamp 1626908933
transform 1 0 29184 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_47
timestamp 1626908933
transform 1 0 29184 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1394
timestamp 1626908933
transform 1 0 29568 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_403
timestamp 1626908933
transform 1 0 29568 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_797
timestamp 1626908933
transform 1 0 29664 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_75
timestamp 1626908933
transform 1 0 29664 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1393
timestamp 1626908933
transform 1 0 30432 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_402
timestamp 1626908933
transform 1 0 30432 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_619
timestamp 1626908933
transform 1 0 30528 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_21
timestamp 1626908933
transform 1 0 30528 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_751
timestamp 1626908933
transform 1 0 30912 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_29
timestamp 1626908933
transform 1 0 30912 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_224
timestamp 1626908933
transform 1 0 31680 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_581
timestamp 1626908933
transform 1 0 31680 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_445
timestamp 1626908933
transform 1 0 31776 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1046
timestamp 1626908933
transform 1 0 31776 0 -1 11988
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_15
timestamp 1626908933
transform 1 0 31700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_663
timestamp 1626908933
transform 1 0 31700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_15
timestamp 1626908933
transform 1 0 31700 0 1 11322
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_663
timestamp 1626908933
transform 1 0 31700 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_797
timestamp 1626908933
transform 1 0 31968 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1788
timestamp 1626908933
transform 1 0 31968 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3875
timestamp 1626908933
transform 1 0 144 0 1 11507
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1908
timestamp 1626908933
transform 1 0 144 0 1 11507
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1789
timestamp 1626908933
transform 1 0 192 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_798
timestamp 1626908933
transform 1 0 192 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1790
timestamp 1626908933
transform 1 0 384 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_799
timestamp 1626908933
transform 1 0 384 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_580
timestamp 1626908933
transform 1 0 288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_223
timestamp 1626908933
transform 1 0 288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1047
timestamp 1626908933
transform 1 0 0 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_446
timestamp 1626908933
transform 1 0 0 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1
timestamp 1626908933
transform 1 0 624 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1968
timestamp 1626908933
transform 1 0 624 0 1 11581
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1
timestamp 1626908933
transform 1 0 624 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1875
timestamp 1626908933
transform 1 0 720 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1936
timestamp 1626908933
transform 1 0 624 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3810
timestamp 1626908933
transform 1 0 720 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_3
timestamp 1626908933
transform -1 0 1344 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_11
timestamp 1626908933
transform -1 0 1344 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_447
timestamp 1626908933
transform 1 0 1344 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1048
timestamp 1626908933
transform 1 0 1344 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_7
timestamp 1626908933
transform 1 0 1200 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1317
timestamp 1626908933
transform 1 0 1392 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1974
timestamp 1626908933
transform 1 0 1200 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3284
timestamp 1626908933
transform 1 0 1392 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_9
timestamp 1626908933
transform 1 0 1200 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1944
timestamp 1626908933
transform 1 0 1200 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_800
timestamp 1626908933
transform 1 0 1536 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1791
timestamp 1626908933
transform 1 0 1536 0 1 11988
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_639
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1287
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_639
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1287
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_2
timestamp 1626908933
transform 1 0 1632 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_10
timestamp 1626908933
transform 1 0 1632 0 1 11988
box -38 -49 902 715
use M1M2_PR  M1M2_PR_2276
timestamp 1626908933
transform 1 0 2256 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_309
timestamp 1626908933
transform 1 0 2256 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1792
timestamp 1626908933
transform 1 0 2688 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_801
timestamp 1626908933
transform 1 0 2688 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1049
timestamp 1626908933
transform 1 0 2496 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_448
timestamp 1626908933
transform 1 0 2496 0 1 11988
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1263
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_615
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1263
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_615
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3332
timestamp 1626908933
transform 1 0 3888 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2268
timestamp 1626908933
transform 1 0 2928 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1397
timestamp 1626908933
transform 1 0 3888 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_333
timestamp 1626908933
transform 1 0 2928 0 1 12099
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_519
timestamp 1626908933
transform 1 0 4608 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1117
timestamp 1626908933
transform 1 0 4608 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_401
timestamp 1626908933
transform 1 0 4512 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1392
timestamp 1626908933
transform 1 0 4512 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1474
timestamp 1626908933
transform 1 0 4272 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3409
timestamp 1626908933
transform 1 0 4272 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_222
timestamp 1626908933
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_579
timestamp 1626908933
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1389
timestamp 1626908933
transform 1 0 4848 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3356
timestamp 1626908933
transform 1 0 4848 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_449
timestamp 1626908933
transform 1 0 5376 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1050
timestamp 1626908933
transform 1 0 5376 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_0
timestamp 1626908933
transform 1 0 5088 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_5
timestamp 1626908933
transform 1 0 5088 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_9
timestamp 1626908933
transform -1 0 4512 0 1 11988
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_3
timestamp 1626908933
transform -1 0 4512 0 1 11988
box -38 -49 1766 715
use M1M2_PR  M1M2_PR_1319
timestamp 1626908933
transform 1 0 5808 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3286
timestamp 1626908933
transform 1 0 5808 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1399
timestamp 1626908933
transform 1 0 6192 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3334
timestamp 1626908933
transform 1 0 6192 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1468
timestamp 1626908933
transform 1 0 6576 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3403
timestamp 1626908933
transform 1 0 6576 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_706
timestamp 1626908933
transform 1 0 6864 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2673
timestamp 1626908933
transform 1 0 6864 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_902
timestamp 1626908933
transform 1 0 7056 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2869
timestamp 1626908933
transform 1 0 7056 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_952
timestamp 1626908933
transform 1 0 7056 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2887
timestamp 1626908933
transform 1 0 7056 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_726
timestamp 1626908933
transform 1 0 7248 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2661
timestamp 1626908933
transform 1 0 7248 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_899
timestamp 1626908933
transform 1 0 7344 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2866
timestamp 1626908933
transform 1 0 7344 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_948
timestamp 1626908933
transform 1 0 7344 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2883
timestamp 1626908933
transform 1 0 7344 0 1 11729
box -29 -23 29 23
use M1M2_PR  M1M2_PR_805
timestamp 1626908933
transform 1 0 8112 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2772
timestamp 1626908933
transform 1 0 8112 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_321
timestamp 1626908933
transform 1 0 6192 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2288
timestamp 1626908933
transform 1 0 6192 0 1 12099
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_591
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1239
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_591
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1239
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use M1M2_PR  M1M2_PR_705
timestamp 1626908933
transform 1 0 6864 0 1 12173
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2672
timestamp 1626908933
transform 1 0 6864 0 1 12173
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1531
timestamp 1626908933
transform 1 0 7152 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3498
timestamp 1626908933
transform 1 0 7152 0 1 11877
box -32 -32 32 32
use L1M1_PR  L1M1_PR_347
timestamp 1626908933
transform 1 0 7152 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1618
timestamp 1626908933
transform 1 0 7152 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2282
timestamp 1626908933
transform 1 0 7152 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3553
timestamp 1626908933
transform 1 0 7152 0 1 11877
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_34
timestamp 1626908933
transform -1 0 9504 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_9
timestamp 1626908933
transform -1 0 9504 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_7
timestamp 1626908933
transform 1 0 5568 0 1 11988
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_1
timestamp 1626908933
transform 1 0 5568 0 1 11988
box -38 -49 1766 715
use L1M1_PR  L1M1_PR_839
timestamp 1626908933
transform 1 0 8688 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2774
timestamp 1626908933
transform 1 0 8688 0 1 11581
box -29 -23 29 23
use M1M2_PR  M1M2_PR_802
timestamp 1626908933
transform 1 0 8880 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2769
timestamp 1626908933
transform 1 0 8880 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_836
timestamp 1626908933
transform 1 0 8880 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2771
timestamp 1626908933
transform 1 0 8880 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_808
timestamp 1626908933
transform 1 0 9072 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2775
timestamp 1626908933
transform 1 0 9072 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_842
timestamp 1626908933
transform 1 0 9072 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2777
timestamp 1626908933
transform 1 0 9072 0 1 11729
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_567
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1215
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_567
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1215
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2660
timestamp 1626908933
transform 1 0 9648 0 1 12173
box -29 -23 29 23
use L1M1_PR  L1M1_PR_725
timestamp 1626908933
transform 1 0 9648 0 1 12173
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2670
timestamp 1626908933
transform 1 0 9648 0 1 12173
box -32 -32 32 32
use M1M2_PR  M1M2_PR_703
timestamp 1626908933
transform 1 0 9648 0 1 12173
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_578
timestamp 1626908933
transform 1 0 9984 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_221
timestamp 1626908933
transform 1 0 9984 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_28
timestamp 1626908933
transform 1 0 9504 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_97
timestamp 1626908933
transform 1 0 9504 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_209
timestamp 1626908933
transform 1 0 10080 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_810
timestamp 1626908933
transform 1 0 10080 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_2923
timestamp 1626908933
transform 1 0 10608 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_988
timestamp 1626908933
transform 1 0 10608 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2901
timestamp 1626908933
transform 1 0 10608 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_934
timestamp 1626908933
transform 1 0 10608 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2920
timestamp 1626908933
transform 1 0 10800 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_985
timestamp 1626908933
transform 1 0 10800 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3534
timestamp 1626908933
transform 1 0 10416 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1599
timestamp 1626908933
transform 1 0 10416 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3480
timestamp 1626908933
transform 1 0 10416 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1513
timestamp 1626908933
transform 1 0 10416 0 1 11877
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_517
timestamp 1626908933
transform 1 0 10272 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1239
timestamp 1626908933
transform 1 0 10272 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2095
timestamp 1626908933
transform 1 0 10896 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_160
timestamp 1626908933
transform 1 0 10896 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2111
timestamp 1626908933
transform 1 0 10896 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_144
timestamp 1626908933
transform 1 0 10896 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_91
timestamp 1626908933
transform 1 0 11040 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_30
timestamp 1626908933
transform 1 0 11040 0 1 11988
box -38 -49 326 715
use M1M2_PR  M1M2_PR_770
timestamp 1626908933
transform 1 0 11568 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2737
timestamp 1626908933
transform 1 0 11568 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_931
timestamp 1626908933
transform 1 0 11088 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2898
timestamp 1626908933
transform 1 0 11088 0 1 11877
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_543
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1191
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_543
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1191
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_75
timestamp 1626908933
transform -1 0 12192 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_6
timestamp 1626908933
transform -1 0 12192 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_27
timestamp 1626908933
transform 1 0 11328 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_79
timestamp 1626908933
transform 1 0 11328 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_208
timestamp 1626908933
transform 1 0 12192 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_809
timestamp 1626908933
transform 1 0 12192 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_151
timestamp 1626908933
transform 1 0 12144 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_152
timestamp 1626908933
transform 1 0 12048 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2118
timestamp 1626908933
transform 1 0 12144 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2119
timestamp 1626908933
transform 1 0 12048 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_400
timestamp 1626908933
transform 1 0 12384 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1391
timestamp 1626908933
transform 1 0 12384 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_371
timestamp 1626908933
transform 1 0 12480 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_969
timestamp 1626908933
transform 1 0 12480 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_207
timestamp 1626908933
transform 1 0 13440 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_808
timestamp 1626908933
transform 1 0 13440 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_672
timestamp 1626908933
transform 1 0 13200 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2639
timestamp 1626908933
transform 1 0 13200 0 1 11581
box -32 -32 32 32
use L1M1_PR  L1M1_PR_168
timestamp 1626908933
transform 1 0 13392 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_689
timestamp 1626908933
transform 1 0 13488 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2103
timestamp 1626908933
transform 1 0 13392 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2624
timestamp 1626908933
transform 1 0 13488 0 1 11581
box -29 -23 29 23
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_2
timestamp 1626908933
transform -1 0 13440 0 1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_6
timestamp 1626908933
transform -1 0 13440 0 1 11988
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1167
timestamp 1626908933
transform 1 0 13700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_519
timestamp 1626908933
transform 1 0 13700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1167
timestamp 1626908933
transform 1 0 13700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_519
timestamp 1626908933
transform 1 0 13700 0 1 11988
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2735
timestamp 1626908933
transform 1 0 13776 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_768
timestamp 1626908933
transform 1 0 13776 0 1 11803
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1165
timestamp 1626908933
transform 1 0 13632 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_443
timestamp 1626908933
transform 1 0 13632 0 1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_54
timestamp 1626908933
transform 1 0 14064 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2021
timestamp 1626908933
transform 1 0 14064 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1666
timestamp 1626908933
transform 1 0 14256 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3633
timestamp 1626908933
transform 1 0 14256 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_61
timestamp 1626908933
transform 1 0 13872 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_800
timestamp 1626908933
transform 1 0 13968 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1996
timestamp 1626908933
transform 1 0 13872 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2735
timestamp 1626908933
transform 1 0 13968 0 1 11729
box -29 -23 29 23
use M1M2_PR  M1M2_PR_150
timestamp 1626908933
transform 1 0 13872 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2117
timestamp 1626908933
transform 1 0 13872 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_64
timestamp 1626908933
transform -1 0 14688 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_2
timestamp 1626908933
transform -1 0 14688 0 1 11988
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2100
timestamp 1626908933
transform 1 0 14736 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_165
timestamp 1626908933
transform 1 0 14736 0 1 12099
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1793
timestamp 1626908933
transform 1 0 14880 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_802
timestamp 1626908933
transform 1 0 14880 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1051
timestamp 1626908933
transform 1 0 14688 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_450
timestamp 1626908933
transform 1 0 14688 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1052
timestamp 1626908933
transform 1 0 15456 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_451
timestamp 1626908933
transform 1 0 15456 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_919
timestamp 1626908933
transform 1 0 15072 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_321
timestamp 1626908933
transform 1 0 15072 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_577
timestamp 1626908933
transform 1 0 14976 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_220
timestamp 1626908933
transform 1 0 14976 0 1 11988
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1143
timestamp 1626908933
transform 1 0 16100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_495
timestamp 1626908933
transform 1 0 16100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1143
timestamp 1626908933
transform 1 0 16100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_495
timestamp 1626908933
transform 1 0 16100 0 1 11988
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3678
timestamp 1626908933
transform 1 0 15504 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1711
timestamp 1626908933
transform 1 0 15504 0 1 11581
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_20
timestamp 1626908933
transform 1 0 15648 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_89
timestamp 1626908933
transform 1 0 15648 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1053
timestamp 1626908933
transform 1 0 16512 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_452
timestamp 1626908933
transform 1 0 16512 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_900
timestamp 1626908933
transform 1 0 16128 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_302
timestamp 1626908933
transform 1 0 16128 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_85
timestamp 1626908933
transform -1 0 16992 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_23
timestamp 1626908933
transform -1 0 16992 0 1 11988
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3682
timestamp 1626908933
transform 1 0 16752 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1747
timestamp 1626908933
transform 1 0 16752 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3434
timestamp 1626908933
transform 1 0 16944 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1467
timestamp 1626908933
transform 1 0 16944 0 1 11729
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_80
timestamp 1626908933
transform 1 0 16992 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_28
timestamp 1626908933
transform 1 0 16992 0 1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3486
timestamp 1626908933
transform 1 0 17136 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1551
timestamp 1626908933
transform 1 0 17136 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1054
timestamp 1626908933
transform 1 0 17376 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_453
timestamp 1626908933
transform 1 0 17376 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_77
timestamp 1626908933
transform 1 0 17568 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_15
timestamp 1626908933
transform 1 0 17568 0 1 11988
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2751
timestamp 1626908933
transform 1 0 17712 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_816
timestamp 1626908933
transform 1 0 17712 0 1 12099
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_807
timestamp 1626908933
transform 1 0 17856 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_206
timestamp 1626908933
transform 1 0 17856 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_2751
timestamp 1626908933
transform 1 0 18000 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2551
timestamp 1626908933
transform 1 0 18096 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_784
timestamp 1626908933
transform 1 0 18000 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_584
timestamp 1626908933
transform 1 0 18096 0 1 11581
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1794
timestamp 1626908933
transform 1 0 18432 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_803
timestamp 1626908933
transform 1 0 18432 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_849
timestamp 1626908933
transform 1 0 18048 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_251
timestamp 1626908933
transform 1 0 18048 0 1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_695
timestamp 1626908933
transform 1 0 18768 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2630
timestamp 1626908933
transform 1 0 18768 0 1 12099
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_471
timestamp 1626908933
transform 1 0 18500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1119
timestamp 1626908933
transform 1 0 18500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_471
timestamp 1626908933
transform 1 0 18500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1119
timestamp 1626908933
transform 1 0 18500 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_3
timestamp 1626908933
transform 1 0 18528 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_64
timestamp 1626908933
transform 1 0 18528 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_245
timestamp 1626908933
transform 1 0 18816 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_843
timestamp 1626908933
transform 1 0 18816 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2644
timestamp 1626908933
transform 1 0 19056 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_677
timestamp 1626908933
transform 1 0 19056 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1055
timestamp 1626908933
transform 1 0 19200 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_454
timestamp 1626908933
transform 1 0 19200 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_455
timestamp 1626908933
transform 1 0 19680 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1056
timestamp 1626908933
transform 1 0 19680 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_697
timestamp 1626908933
transform 1 0 19536 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2632
timestamp 1626908933
transform 1 0 19536 0 1 12099
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_219
timestamp 1626908933
transform 1 0 19968 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_576
timestamp 1626908933
transform 1 0 19968 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_804
timestamp 1626908933
transform 1 0 19872 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1795
timestamp 1626908933
transform 1 0 19872 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_678
timestamp 1626908933
transform 1 0 19920 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2645
timestamp 1626908933
transform 1 0 19920 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_11
timestamp 1626908933
transform -1 0 19680 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_73
timestamp 1626908933
transform -1 0 19680 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_46
timestamp 1626908933
transform -1 0 21216 0 1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_7
timestamp 1626908933
transform -1 0 21216 0 1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_806
timestamp 1626908933
transform 1 0 20064 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_205
timestamp 1626908933
transform 1 0 20064 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_815
timestamp 1626908933
transform 1 0 20256 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_217
timestamp 1626908933
transform 1 0 20256 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_77
timestamp 1626908933
transform 1 0 20688 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2044
timestamp 1626908933
transform 1 0 20688 0 1 11729
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_447
timestamp 1626908933
transform 1 0 20900 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1095
timestamp 1626908933
transform 1 0 20900 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_447
timestamp 1626908933
transform 1 0 20900 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1095
timestamp 1626908933
transform 1 0 20900 0 1 11988
box -100 -49 100 49
use M1M2_PR  M1M2_PR_866
timestamp 1626908933
transform 1 0 21072 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2833
timestamp 1626908933
transform 1 0 21072 0 1 11877
box -32 -32 32 32
use L1M1_PR  L1M1_PR_85
timestamp 1626908933
transform 1 0 21072 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_912
timestamp 1626908933
transform 1 0 21072 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2020
timestamp 1626908933
transform 1 0 21072 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2847
timestamp 1626908933
transform 1 0 21072 0 1 11877
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_204
timestamp 1626908933
transform 1 0 21216 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_805
timestamp 1626908933
transform 1 0 21216 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_864
timestamp 1626908933
transform 1 0 21264 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2831
timestamp 1626908933
transform 1 0 21264 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_907
timestamp 1626908933
transform 1 0 21264 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2842
timestamp 1626908933
transform 1 0 21264 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_805
timestamp 1626908933
transform 1 0 21792 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1796
timestamp 1626908933
transform 1 0 21792 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_789
timestamp 1626908933
transform 1 0 21936 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2756
timestamp 1626908933
transform 1 0 21936 0 1 11803
box -32 -32 32 32
use L1M1_PR  L1M1_PR_590
timestamp 1626908933
transform 1 0 21936 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2525
timestamp 1626908933
transform 1 0 21936 0 1 11581
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_196
timestamp 1626908933
transform 1 0 21408 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_794
timestamp 1626908933
transform 1 0 21408 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_19
timestamp 1626908933
transform -1 0 22176 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_81
timestamp 1626908933
transform -1 0 22176 0 1 11988
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2852
timestamp 1626908933
transform 1 0 22032 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2489
timestamp 1626908933
transform 1 0 22032 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_917
timestamp 1626908933
transform 1 0 22032 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_554
timestamp 1626908933
transform 1 0 22032 0 1 11729
box -29 -23 29 23
use M1M2_PR  M1M2_PR_788
timestamp 1626908933
transform 1 0 22320 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2755
timestamp 1626908933
transform 1 0 22320 0 1 11581
box -32 -32 32 32
use L1M1_PR  L1M1_PR_819
timestamp 1626908933
transform 1 0 22320 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2754
timestamp 1626908933
transform 1 0 22320 0 1 11581
box -29 -23 29 23
use M1M2_PR  M1M2_PR_166
timestamp 1626908933
transform 1 0 22416 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2133
timestamp 1626908933
transform 1 0 22416 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_183
timestamp 1626908933
transform 1 0 22416 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2118
timestamp 1626908933
transform 1 0 22416 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_547
timestamp 1626908933
transform 1 0 22512 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2514
timestamp 1626908933
transform 1 0 22512 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_821
timestamp 1626908933
transform 1 0 22128 0 1 11803
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2756
timestamp 1626908933
transform 1 0 22128 0 1 11803
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_804
timestamp 1626908933
transform 1 0 22176 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_203
timestamp 1626908933
transform 1 0 22176 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_177
timestamp 1626908933
transform 1 0 22368 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_775
timestamp 1626908933
transform 1 0 22368 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_21
timestamp 1626908933
transform 1 0 22752 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_83
timestamp 1626908933
transform 1 0 22752 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_399
timestamp 1626908933
transform 1 0 23136 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1390
timestamp 1626908933
transform 1 0 23136 0 1 11988
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_423
timestamp 1626908933
transform 1 0 23300 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1071
timestamp 1626908933
transform 1 0 23300 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_423
timestamp 1626908933
transform 1 0 23300 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1071
timestamp 1626908933
transform 1 0 23300 0 1 11988
box -100 -49 100 49
use M1M2_PR  M1M2_PR_565
timestamp 1626908933
transform 1 0 23760 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_869
timestamp 1626908933
transform 1 0 23568 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_870
timestamp 1626908933
transform 1 0 23568 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2532
timestamp 1626908933
transform 1 0 23760 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2836
timestamp 1626908933
transform 1 0 23568 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2837
timestamp 1626908933
transform 1 0 23568 0 1 11877
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_234
timestamp 1626908933
transform 1 0 23232 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_956
timestamp 1626908933
transform 1 0 23232 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2504
timestamp 1626908933
transform 1 0 24240 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_569
timestamp 1626908933
transform 1 0 24240 0 1 12099
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1389
timestamp 1626908933
transform 1 0 24288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_398
timestamp 1626908933
transform 1 0 24288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_741
timestamp 1626908933
transform 1 0 24384 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_143
timestamp 1626908933
transform 1 0 24384 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_66
timestamp 1626908933
transform 1 0 24000 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_5
timestamp 1626908933
transform 1 0 24000 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1797
timestamp 1626908933
transform 1 0 24864 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1388
timestamp 1626908933
transform 1 0 24768 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_806
timestamp 1626908933
transform 1 0 24864 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_397
timestamp 1626908933
transform 1 0 24768 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_218
timestamp 1626908933
transform 1 0 24960 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_575
timestamp 1626908933
transform 1 0 24960 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_396
timestamp 1626908933
transform 1 0 25056 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1387
timestamp 1626908933
transform 1 0 25056 0 1 11988
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_399
timestamp 1626908933
transform 1 0 25700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1047
timestamp 1626908933
transform 1 0 25700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_399
timestamp 1626908933
transform 1 0 25700 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1047
timestamp 1626908933
transform 1 0 25700 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_124
timestamp 1626908933
transform 1 0 25152 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_722
timestamp 1626908933
transform 1 0 25152 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_34
timestamp 1626908933
transform 1 0 25536 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_96
timestamp 1626908933
transform 1 0 25536 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1386
timestamp 1626908933
transform 1 0 25920 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_395
timestamp 1626908933
transform 1 0 25920 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_881
timestamp 1626908933
transform 1 0 26016 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_159
timestamp 1626908933
transform 1 0 26016 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2033
timestamp 1626908933
transform 1 0 27312 0 1 12173
box -29 -23 29 23
use L1M1_PR  L1M1_PR_98
timestamp 1626908933
transform 1 0 27312 0 1 12173
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1385
timestamp 1626908933
transform 1 0 27264 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_394
timestamp 1626908933
transform 1 0 27264 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_683
timestamp 1626908933
transform 1 0 27360 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_85
timestamp 1626908933
transform 1 0 27360 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_4
timestamp 1626908933
transform -1 0 27264 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_73
timestamp 1626908933
transform -1 0 27264 0 1 11988
box -38 -49 518 715
use L1M1_PR  L1M1_PR_97
timestamp 1626908933
transform 1 0 28176 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2032
timestamp 1626908933
transform 1 0 28176 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_915
timestamp 1626908933
transform 1 0 27888 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2850
timestamp 1626908933
transform 1 0 27888 0 1 11877
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_375
timestamp 1626908933
transform 1 0 28100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1023
timestamp 1626908933
transform 1 0 28100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_375
timestamp 1626908933
transform 1 0 28100 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1023
timestamp 1626908933
transform 1 0 28100 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_127
timestamp 1626908933
transform 1 0 27744 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_849
timestamp 1626908933
transform 1 0 27744 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_202
timestamp 1626908933
transform 1 0 28512 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_803
timestamp 1626908933
transform 1 0 28512 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_393
timestamp 1626908933
transform 1 0 28704 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1384
timestamp 1626908933
transform 1 0 28704 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_86
timestamp 1626908933
transform 1 0 28560 0 1 12173
box -32 -32 32 32
use M1M2_PR  M1M2_PR_87
timestamp 1626908933
transform 1 0 28560 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2053
timestamp 1626908933
transform 1 0 28560 0 1 12173
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2054
timestamp 1626908933
transform 1 0 28560 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_868
timestamp 1626908933
transform 1 0 28944 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2835
timestamp 1626908933
transform 1 0 28944 0 1 11877
box -32 -32 32 32
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_8
timestamp 1626908933
transform 1 0 28800 0 1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_47
timestamp 1626908933
transform 1 0 28800 0 1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_201
timestamp 1626908933
transform 1 0 29376 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_802
timestamp 1626908933
transform 1 0 29376 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_96
timestamp 1626908933
transform 1 0 29424 0 1 12173
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2031
timestamp 1626908933
transform 1 0 29424 0 1 12173
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_217
timestamp 1626908933
transform 1 0 29952 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_574
timestamp 1626908933
transform 1 0 29952 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_200
timestamp 1626908933
transform 1 0 30048 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_801
timestamp 1626908933
transform 1 0 30048 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_44
timestamp 1626908933
transform 1 0 29568 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_642
timestamp 1626908933
transform 1 0 29568 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1383
timestamp 1626908933
transform 1 0 30240 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_392
timestamp 1626908933
transform 1 0 30240 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_773
timestamp 1626908933
transform 1 0 30336 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_51
timestamp 1626908933
transform 1 0 30336 0 1 11988
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_999
timestamp 1626908933
transform 1 0 30500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_351
timestamp 1626908933
transform 1 0 30500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_999
timestamp 1626908933
transform 1 0 30500 0 1 11988
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_351
timestamp 1626908933
transform 1 0 30500 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1382
timestamp 1626908933
transform 1 0 31104 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_391
timestamp 1626908933
transform 1 0 31104 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_736
timestamp 1626908933
transform 1 0 31200 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_14
timestamp 1626908933
transform 1 0 31200 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1798
timestamp 1626908933
transform 1 0 31968 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_807
timestamp 1626908933
transform 1 0 31968 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_199
timestamp 1626908933
transform 1 0 0 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_800
timestamp 1626908933
transform 1 0 0 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1907
timestamp 1626908933
transform 1 0 144 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3874
timestamp 1626908933
transform 1 0 144 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_0
timestamp 1626908933
transform 1 0 624 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1967
timestamp 1626908933
transform 1 0 624 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_0
timestamp 1626908933
transform 1 0 624 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1935
timestamp 1626908933
transform 1 0 624 0 1 12321
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_326
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_974
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_326
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_974
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_714
timestamp 1626908933
transform 1 0 192 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1436
timestamp 1626908933
transform 1 0 192 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_390
timestamp 1626908933
transform 1 0 960 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1381
timestamp 1626908933
transform 1 0 960 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_7
timestamp 1626908933
transform 1 0 1200 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1873
timestamp 1626908933
transform 1 0 912 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1942
timestamp 1626908933
transform 1 0 1200 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3808
timestamp 1626908933
transform 1 0 912 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_5
timestamp 1626908933
transform 1 0 1488 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1906
timestamp 1626908933
transform 1 0 1392 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1972
timestamp 1626908933
transform 1 0 1488 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3873
timestamp 1626908933
transform 1 0 1392 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_680
timestamp 1626908933
transform 1 0 1440 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1402
timestamp 1626908933
transform 1 0 1440 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_576
timestamp 1626908933
transform 1 0 1056 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1174
timestamp 1626908933
transform 1 0 1056 0 -1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_4
timestamp 1626908933
transform 1 0 1776 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1870
timestamp 1626908933
transform 1 0 1776 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1939
timestamp 1626908933
transform 1 0 1776 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3805
timestamp 1626908933
transform 1 0 1776 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_389
timestamp 1626908933
transform 1 0 2208 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1380
timestamp 1626908933
transform 1 0 2208 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_6
timestamp 1626908933
transform 1 0 2160 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1941
timestamp 1626908933
transform 1 0 2160 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_216
timestamp 1626908933
transform 1 0 2496 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_573
timestamp 1626908933
transform 1 0 2496 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_456
timestamp 1626908933
transform 1 0 2304 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1057
timestamp 1626908933
transform 1 0 2304 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1965
timestamp 1626908933
transform 1 0 2448 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3932
timestamp 1626908933
transform 1 0 2448 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1379
timestamp 1626908933
transform 1 0 2592 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_388
timestamp 1626908933
transform 1 0 2592 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1377
timestamp 1626908933
transform 1 0 2688 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_655
timestamp 1626908933
transform 1 0 2688 0 -1 13320
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_302
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_950
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_302
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_950
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_3
timestamp 1626908933
transform 1 0 3456 0 -1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_1
timestamp 1626908933
transform 1 0 3456 0 -1 13320
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1393
timestamp 1626908933
transform 1 0 3696 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3360
timestamp 1626908933
transform 1 0 3696 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1315
timestamp 1626908933
transform 1 0 3888 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3282
timestamp 1626908933
transform 1 0 3888 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1395
timestamp 1626908933
transform 1 0 4080 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1475
timestamp 1626908933
transform 1 0 3984 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3330
timestamp 1626908933
transform 1 0 4080 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3410
timestamp 1626908933
transform 1 0 3984 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1473
timestamp 1626908933
transform 1 0 4560 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3408
timestamp 1626908933
transform 1 0 4560 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1321
timestamp 1626908933
transform 1 0 5040 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1388
timestamp 1626908933
transform 1 0 4848 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3288
timestamp 1626908933
transform 1 0 5040 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3355
timestamp 1626908933
transform 1 0 4848 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1402
timestamp 1626908933
transform 1 0 5136 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3337
timestamp 1626908933
transform 1 0 5136 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_429
timestamp 1626908933
transform 1 0 5232 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2364
timestamp 1626908933
transform 1 0 5232 0 1 12543
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_278
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_926
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_278
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_926
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1387
timestamp 1626908933
transform 1 0 4848 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3354
timestamp 1626908933
transform 1 0 4848 0 1 12765
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1470
timestamp 1626908933
transform 1 0 5232 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3405
timestamp 1626908933
transform 1 0 5232 0 1 12765
box -29 -23 29 23
use M1M2_PR  M1M2_PR_428
timestamp 1626908933
transform 1 0 5520 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2395
timestamp 1626908933
transform 1 0 5520 0 1 12765
box -32 -32 32 32
use sky130_fd_sc_hs__sdlclkp_1  sky130_fd_sc_hs__sdlclkp_1_1
timestamp 1626908933
transform 1 0 3744 0 -1 13320
box -38 -49 1574 715
use sky130_fd_sc_hs__sdlclkp_1  sky130_fd_sc_hs__sdlclkp_1_0
timestamp 1626908933
transform 1 0 3744 0 -1 13320
box -38 -49 1574 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_6
timestamp 1626908933
transform 1 0 5280 0 -1 13320
box -38 -49 1766 715
use sky130_fd_sc_hs__dfxtp_2  sky130_fd_sc_hs__dfxtp_2_0
timestamp 1626908933
transform 1 0 5280 0 -1 13320
box -38 -49 1766 715
use L1M1_PR  L1M1_PR_3404
timestamp 1626908933
transform 1 0 5616 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3336
timestamp 1626908933
transform 1 0 6000 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2357
timestamp 1626908933
transform 1 0 6864 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1469
timestamp 1626908933
transform 1 0 5616 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1401
timestamp 1626908933
transform 1 0 6000 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_422
timestamp 1626908933
transform 1 0 6864 0 1 12765
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2400
timestamp 1626908933
transform 1 0 5808 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_433
timestamp 1626908933
transform 1 0 5808 0 1 12543
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_475
timestamp 1626908933
transform 1 0 7104 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1073
timestamp 1626908933
transform 1 0 7104 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_387
timestamp 1626908933
transform 1 0 7008 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1378
timestamp 1626908933
transform 1 0 7008 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1530
timestamp 1626908933
transform 1 0 7152 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3497
timestamp 1626908933
transform 1 0 7152 0 1 12913
box -32 -32 32 32
use L1M1_PR  L1M1_PR_161
timestamp 1626908933
transform 1 0 7344 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2096
timestamp 1626908933
transform 1 0 7344 0 1 12469
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_215
timestamp 1626908933
transform 1 0 7488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_572
timestamp 1626908933
transform 1 0 7488 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1617
timestamp 1626908933
transform 1 0 7632 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3552
timestamp 1626908933
transform 1 0 7632 0 1 12913
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_254
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_902
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_254
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_902
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1672
timestamp 1626908933
transform 1 0 8016 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3639
timestamp 1626908933
transform 1 0 8016 0 1 12247
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_25
timestamp 1626908933
transform 1 0 7584 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_0
timestamp 1626908933
transform 1 0 7584 0 -1 13320
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_3688
timestamp 1626908933
transform 1 0 9168 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3535
timestamp 1626908933
transform 1 0 9456 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1753
timestamp 1626908933
transform 1 0 9168 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1600
timestamp 1626908933
transform 1 0 9456 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3706
timestamp 1626908933
transform 1 0 8304 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3705
timestamp 1626908933
transform 1 0 8304 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1739
timestamp 1626908933
transform 1 0 8304 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1738
timestamp 1626908933
transform 1 0 8304 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2065
timestamp 1626908933
transform 1 0 9744 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_130
timestamp 1626908933
transform 1 0 9744 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2086
timestamp 1626908933
transform 1 0 9744 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_119
timestamp 1626908933
transform 1 0 9744 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2064
timestamp 1626908933
transform 1 0 9744 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_129
timestamp 1626908933
transform 1 0 9744 0 1 12765
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2085
timestamp 1626908933
transform 1 0 9744 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_118
timestamp 1626908933
transform 1 0 9744 0 1 12765
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1799
timestamp 1626908933
transform 1 0 9792 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_808
timestamp 1626908933
transform 1 0 9792 0 -1 13320
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_230
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_878
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_230
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_878
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use M1M2_PR  M1M2_PR_147
timestamp 1626908933
transform 1 0 10416 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_661
timestamp 1626908933
transform 1 0 10320 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1512
timestamp 1626908933
transform 1 0 10416 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2114
timestamp 1626908933
transform 1 0 10416 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2628
timestamp 1626908933
transform 1 0 10320 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3479
timestamp 1626908933
transform 1 0 10416 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_933
timestamp 1626908933
transform 1 0 10608 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2900
timestamp 1626908933
transform 1 0 10608 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_143
timestamp 1626908933
transform 1 0 10896 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2110
timestamp 1626908933
transform 1 0 10896 0 1 12469
box -32 -32 32 32
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_34
timestamp 1626908933
transform 1 0 9888 0 -1 13320
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_10
timestamp 1626908933
transform 1 0 9888 0 -1 13320
box -38 -49 2342 715
use L1M1_PR  L1M1_PR_2921
timestamp 1626908933
transform 1 0 11184 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2919
timestamp 1626908933
transform 1 0 11088 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2093
timestamp 1626908933
transform 1 0 11376 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_986
timestamp 1626908933
transform 1 0 11184 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_984
timestamp 1626908933
transform 1 0 11088 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_158
timestamp 1626908933
transform 1 0 11376 0 1 12469
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2897
timestamp 1626908933
transform 1 0 11088 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_930
timestamp 1626908933
transform 1 0 11088 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2625
timestamp 1626908933
transform 1 0 12048 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2004
timestamp 1626908933
transform 1 0 11856 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2000
timestamp 1626908933
transform 1 0 12144 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_690
timestamp 1626908933
transform 1 0 12048 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_69
timestamp 1626908933
transform 1 0 11856 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_65
timestamp 1626908933
transform 1 0 12144 0 1 12913
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2029
timestamp 1626908933
transform 1 0 11760 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_62
timestamp 1626908933
transform 1 0 11760 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2624
timestamp 1626908933
transform 1 0 12336 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_657
timestamp 1626908933
transform 1 0 12336 0 1 12395
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_854
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_206
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_854
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_206
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1800
timestamp 1626908933
transform 1 0 12384 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_809
timestamp 1626908933
transform 1 0 12384 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1058
timestamp 1626908933
transform 1 0 12192 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_457
timestamp 1626908933
transform 1 0 12192 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_214
timestamp 1626908933
transform 1 0 12480 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_571
timestamp 1626908933
transform 1 0 12480 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_458
timestamp 1626908933
transform 1 0 12576 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1059
timestamp 1626908933
transform 1 0 12576 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_57
timestamp 1626908933
transform 1 0 12720 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2024
timestamp 1626908933
transform 1 0 12720 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2023
timestamp 1626908933
transform 1 0 12816 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_56
timestamp 1626908933
transform 1 0 12816 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2612
timestamp 1626908933
transform 1 0 12912 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_677
timestamp 1626908933
transform 1 0 12912 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2629
timestamp 1626908933
transform 1 0 12912 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_662
timestamp 1626908933
transform 1 0 12912 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2606
timestamp 1626908933
transform 1 0 13008 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_671
timestamp 1626908933
transform 1 0 13008 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2589
timestamp 1626908933
transform 1 0 13104 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_654
timestamp 1626908933
transform 1 0 13104 0 1 12469
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2638
timestamp 1626908933
transform 1 0 13200 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_671
timestamp 1626908933
transform 1 0 13200 0 1 12543
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_90
timestamp 1626908933
transform -1 0 13248 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_21
timestamp 1626908933
transform -1 0 13248 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_29
timestamp 1626908933
transform 1 0 13248 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_81
timestamp 1626908933
transform 1 0 13248 0 -1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2605
timestamp 1626908933
transform 1 0 13296 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1997
timestamp 1626908933
transform 1 0 13392 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_670
timestamp 1626908933
transform 1 0 13296 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_62
timestamp 1626908933
transform 1 0 13392 0 1 12247
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1801
timestamp 1626908933
transform 1 0 13824 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_810
timestamp 1626908933
transform 1 0 13824 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1060
timestamp 1626908933
transform 1 0 13632 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_459
timestamp 1626908933
transform 1 0 13632 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_386
timestamp 1626908933
transform 1 0 14208 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1377
timestamp 1626908933
transform 1 0 14208 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_53
timestamp 1626908933
transform 1 0 14160 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2020
timestamp 1626908933
transform 1 0 14160 0 1 12913
box -32 -32 32 32
use L1M1_PR  L1M1_PR_810
timestamp 1626908933
transform 1 0 14064 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2745
timestamp 1626908933
transform 1 0 14064 0 1 12765
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_13
timestamp 1626908933
transform -1 0 14208 0 -1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_75
timestamp 1626908933
transform -1 0 14208 0 -1 13320
box -38 -49 326 715
use M1M2_PR  M1M2_PR_778
timestamp 1626908933
transform 1 0 14544 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2745
timestamp 1626908933
transform 1 0 14544 0 1 12765
box -32 -32 32 32
use L1M1_PR  L1M1_PR_162
timestamp 1626908933
transform 1 0 14256 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_669
timestamp 1626908933
transform 1 0 14448 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_688
timestamp 1626908933
transform 1 0 14352 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2097
timestamp 1626908933
transform 1 0 14256 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2604
timestamp 1626908933
transform 1 0 14448 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2623
timestamp 1626908933
transform 1 0 14352 0 1 12543
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_430
timestamp 1626908933
transform 1 0 14304 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1152
timestamp 1626908933
transform 1 0 14304 0 -1 13320
box -38 -49 806 715
use M1M2_PR  M1M2_PR_48
timestamp 1626908933
transform 1 0 14832 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2015
timestamp 1626908933
transform 1 0 14832 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_57
timestamp 1626908933
transform 1 0 15024 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1992
timestamp 1626908933
transform 1 0 15024 0 1 12913
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_182
timestamp 1626908933
transform 1 0 14900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_830
timestamp 1626908933
transform 1 0 14900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_182
timestamp 1626908933
transform 1 0 14900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_830
timestamp 1626908933
transform 1 0 14900 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_18
timestamp 1626908933
transform -1 0 15360 0 -1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_79
timestamp 1626908933
transform -1 0 15360 0 -1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_198
timestamp 1626908933
transform 1 0 15360 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_799
timestamp 1626908933
transform 1 0 15360 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_643
timestamp 1626908933
transform 1 0 15120 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_644
timestamp 1626908933
transform 1 0 15120 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2610
timestamp 1626908933
transform 1 0 15120 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2611
timestamp 1626908933
transform 1 0 15120 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_838
timestamp 1626908933
transform 1 0 15408 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2805
timestamp 1626908933
transform 1 0 15408 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2813
timestamp 1626908933
transform 1 0 15984 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1989
timestamp 1626908933
transform 1 0 15696 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_878
timestamp 1626908933
transform 1 0 15984 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_54
timestamp 1626908933
transform 1 0 15696 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1802
timestamp 1626908933
transform 1 0 16320 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_811
timestamp 1626908933
transform 1 0 16320 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1132
timestamp 1626908933
transform 1 0 15552 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_410
timestamp 1626908933
transform 1 0 15552 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_79
timestamp 1626908933
transform 1 0 16416 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_17
timestamp 1626908933
transform 1 0 16416 0 -1 13320
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2804
timestamp 1626908933
transform 1 0 16560 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2803
timestamp 1626908933
transform 1 0 16560 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2800
timestamp 1626908933
transform 1 0 16464 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_837
timestamp 1626908933
transform 1 0 16560 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_836
timestamp 1626908933
transform 1 0 16560 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_833
timestamp 1626908933
transform 1 0 16464 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3487
timestamp 1626908933
transform 1 0 16752 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2815
timestamp 1626908933
transform 1 0 16752 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2807
timestamp 1626908933
transform 1 0 16752 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1552
timestamp 1626908933
transform 1 0 16752 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_880
timestamp 1626908933
transform 1 0 16752 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_872
timestamp 1626908933
transform 1 0 16752 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1376
timestamp 1626908933
transform 1 0 16800 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_385
timestamp 1626908933
transform 1 0 16800 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3433
timestamp 1626908933
transform 1 0 16944 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1466
timestamp 1626908933
transform 1 0 16944 0 1 12765
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2811
timestamp 1626908933
transform 1 0 17040 0 1 12469
box -29 -23 29 23
use L1M1_PR  L1M1_PR_876
timestamp 1626908933
transform 1 0 17040 0 1 12469
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_806
timestamp 1626908933
transform 1 0 17300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_158
timestamp 1626908933
transform 1 0 17300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_806
timestamp 1626908933
transform 1 0 17300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_158
timestamp 1626908933
transform 1 0 17300 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1803
timestamp 1626908933
transform 1 0 17376 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1375
timestamp 1626908933
transform 1 0 17280 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_812
timestamp 1626908933
transform 1 0 17376 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_384
timestamp 1626908933
transform 1 0 17280 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_288
timestamp 1626908933
transform 1 0 16896 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_886
timestamp 1626908933
transform 1 0 16896 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_213
timestamp 1626908933
transform 1 0 17472 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_570
timestamp 1626908933
transform 1 0 17472 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_592
timestamp 1626908933
transform 1 0 17808 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_663
timestamp 1626908933
transform 1 0 17520 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2527
timestamp 1626908933
transform 1 0 17808 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2598
timestamp 1626908933
transform 1 0 17520 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_583
timestamp 1626908933
transform 1 0 18096 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2550
timestamp 1626908933
transform 1 0 18096 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_357
timestamp 1626908933
transform 1 0 17568 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1079
timestamp 1626908933
transform 1 0 17568 0 -1 13320
box -38 -49 806 715
use M1M2_PR  M1M2_PR_579
timestamp 1626908933
transform 1 0 18288 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_650
timestamp 1626908933
transform 1 0 18480 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2546
timestamp 1626908933
transform 1 0 18288 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2617
timestamp 1626908933
transform 1 0 18480 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_586
timestamp 1626908933
transform 1 0 18480 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_702
timestamp 1626908933
transform 1 0 18576 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2521
timestamp 1626908933
transform 1 0 18480 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2637
timestamp 1626908933
transform 1 0 18576 0 1 12247
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_197
timestamp 1626908933
transform 1 0 19008 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_798
timestamp 1626908933
transform 1 0 19008 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_685
timestamp 1626908933
transform 1 0 19056 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2652
timestamp 1626908933
transform 1 0 19056 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_90
timestamp 1626908933
transform 1 0 18768 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2025
timestamp 1626908933
transform 1 0 18768 0 1 12247
box -29 -23 29 23
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_3
timestamp 1626908933
transform 1 0 18336 0 -1 13320
box -38 -49 710 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_8
timestamp 1626908933
transform 1 0 18336 0 -1 13320
box -38 -49 710 715
use M1M2_PR  M1M2_PR_2047
timestamp 1626908933
transform 1 0 19344 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_80
timestamp 1626908933
transform 1 0 19344 0 1 12247
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1374
timestamp 1626908933
transform 1 0 19200 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_383
timestamp 1626908933
transform 1 0 19200 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1050
timestamp 1626908933
transform 1 0 19296 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_328
timestamp 1626908933
transform 1 0 19296 0 -1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_701
timestamp 1626908933
transform 1 0 19440 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2636
timestamp 1626908933
transform 1 0 19440 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_88
timestamp 1626908933
transform 1 0 19632 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2023
timestamp 1626908933
transform 1 0 19632 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_76
timestamp 1626908933
transform 1 0 20688 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2043
timestamp 1626908933
transform 1 0 20688 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_86
timestamp 1626908933
transform 1 0 20688 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2021
timestamp 1626908933
transform 1 0 20688 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_909
timestamp 1626908933
transform 1 0 20784 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2844
timestamp 1626908933
transform 1 0 20784 0 1 12395
box -29 -23 29 23
use M1M2_PR  M1M2_PR_865
timestamp 1626908933
transform 1 0 21072 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2832
timestamp 1626908933
transform 1 0 21072 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_913
timestamp 1626908933
transform 1 0 20976 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2848
timestamp 1626908933
transform 1 0 20976 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1538
timestamp 1626908933
transform 1 0 21168 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3473
timestamp 1626908933
transform 1 0 21168 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_863
timestamp 1626908933
transform 1 0 21264 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2830
timestamp 1626908933
transform 1 0 21264 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1453
timestamp 1626908933
transform 1 0 21360 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3420
timestamp 1626908933
transform 1 0 21360 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_911
timestamp 1626908933
transform 1 0 21936 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2846
timestamp 1626908933
transform 1 0 21936 0 1 12321
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_134
timestamp 1626908933
transform 1 0 19700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_782
timestamp 1626908933
transform 1 0 19700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_134
timestamp 1626908933
transform 1 0 19700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_782
timestamp 1626908933
transform 1 0 19700 0 1 12654
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1658
timestamp 1626908933
transform 1 0 21552 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3625
timestamp 1626908933
transform 1 0 21552 0 1 12987
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_110
timestamp 1626908933
transform 1 0 22100 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_758
timestamp 1626908933
transform 1 0 22100 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_110
timestamp 1626908933
transform 1 0 22100 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_758
timestamp 1626908933
transform 1 0 22100 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_38
timestamp 1626908933
transform -1 0 22368 0 -1 13320
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_14
timestamp 1626908933
transform -1 0 22368 0 -1 13320
box -38 -49 2342 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_813
timestamp 1626908933
transform 1 0 22368 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1804
timestamp 1626908933
transform 1 0 22368 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_787
timestamp 1626908933
transform 1 0 22320 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2754
timestamp 1626908933
transform 1 0 22320 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_820
timestamp 1626908933
transform 1 0 22128 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2755
timestamp 1626908933
transform 1 0 22128 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_212
timestamp 1626908933
transform 1 0 22464 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_569
timestamp 1626908933
transform 1 0 22464 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_460
timestamp 1626908933
transform 1 0 22560 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1061
timestamp 1626908933
transform 1 0 22560 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_814
timestamp 1626908933
transform 1 0 22752 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1805
timestamp 1626908933
transform 1 0 22752 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_818
timestamp 1626908933
transform 1 0 22896 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_910
timestamp 1626908933
transform 1 0 22800 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1536
timestamp 1626908933
transform 1 0 22896 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2753
timestamp 1626908933
transform 1 0 22896 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2845
timestamp 1626908933
transform 1 0 22800 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3471
timestamp 1626908933
transform 1 0 22896 0 1 12913
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1450
timestamp 1626908933
transform 1 0 22992 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1451
timestamp 1626908933
transform 1 0 22992 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3417
timestamp 1626908933
transform 1 0 22992 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3418
timestamp 1626908933
transform 1 0 22992 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_916
timestamp 1626908933
transform 1 0 23088 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1535
timestamp 1626908933
transform 1 0 23088 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2851
timestamp 1626908933
transform 1 0 23088 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3470
timestamp 1626908933
transform 1 0 23088 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_738
timestamp 1626908933
transform 1 0 23952 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2673
timestamp 1626908933
transform 1 0 23952 0 1 12395
box -29 -23 29 23
use M1M2_PR  M1M2_PR_173
timestamp 1626908933
transform 1 0 24336 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2140
timestamp 1626908933
transform 1 0 24336 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_189
timestamp 1626908933
transform 1 0 24240 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2124
timestamp 1626908933
transform 1 0 24240 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_81
timestamp 1626908933
transform 1 0 24240 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2048
timestamp 1626908933
transform 1 0 24240 0 1 12765
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_86
timestamp 1626908933
transform 1 0 24500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_734
timestamp 1626908933
transform 1 0 24500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_86
timestamp 1626908933
transform 1 0 24500 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_734
timestamp 1626908933
transform 1 0 24500 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_39
timestamp 1626908933
transform 1 0 22848 0 -1 13320
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_15
timestamp 1626908933
transform 1 0 22848 0 -1 13320
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_2681
timestamp 1626908933
transform 1 0 25008 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_714
timestamp 1626908933
transform 1 0 25008 0 1 12395
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2954
timestamp 1626908933
transform 1 0 25584 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1019
timestamp 1626908933
transform 1 0 25584 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2923
timestamp 1626908933
transform 1 0 25488 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_956
timestamp 1626908933
transform 1 0 25488 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2690
timestamp 1626908933
transform 1 0 25680 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_755
timestamp 1626908933
transform 1 0 25680 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2699
timestamp 1626908933
transform 1 0 25680 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_732
timestamp 1626908933
transform 1 0 25680 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_731
timestamp 1626908933
transform 1 0 25680 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2698
timestamp 1626908933
transform 1 0 25680 0 1 12765
box -32 -32 32 32
use L1M1_PR  L1M1_PR_91
timestamp 1626908933
transform 1 0 25104 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2026
timestamp 1626908933
transform 1 0 25104 0 1 12765
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_188
timestamp 1626908933
transform 1 0 25152 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_910
timestamp 1626908933
transform 1 0 25152 0 -1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3517
timestamp 1626908933
transform 1 0 25872 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2958
timestamp 1626908933
transform 1 0 25872 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1582
timestamp 1626908933
transform 1 0 25872 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1023
timestamp 1626908933
transform 1 0 25872 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3462
timestamp 1626908933
transform 1 0 25872 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1495
timestamp 1626908933
transform 1 0 25872 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2695
timestamp 1626908933
transform 1 0 26064 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_728
timestamp 1626908933
transform 1 0 26064 0 1 12765
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1806
timestamp 1626908933
transform 1 0 26112 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_815
timestamp 1626908933
transform 1 0 26112 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1062
timestamp 1626908933
transform 1 0 25920 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_461
timestamp 1626908933
transform 1 0 25920 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_958
timestamp 1626908933
transform 1 0 26256 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1688
timestamp 1626908933
transform 1 0 26448 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2925
timestamp 1626908933
transform 1 0 26256 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3655
timestamp 1626908933
transform 1 0 26448 0 1 12913
box -32 -32 32 32
use L1M1_PR  L1M1_PR_751
timestamp 1626908933
transform 1 0 26352 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2686
timestamp 1626908933
transform 1 0 26352 0 1 12765
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_106
timestamp 1626908933
transform -1 0 26688 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_37
timestamp 1626908933
transform -1 0 26688 0 -1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_736
timestamp 1626908933
transform 1 0 26832 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2671
timestamp 1626908933
transform 1 0 26832 0 1 12395
box -29 -23 29 23
use M1M2_PR  M1M2_PR_176
timestamp 1626908933
transform 1 0 26640 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2143
timestamp 1626908933
transform 1 0 26640 0 1 12987
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_62
timestamp 1626908933
transform 1 0 26900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_710
timestamp 1626908933
transform 1 0 26900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_62
timestamp 1626908933
transform 1 0 26900 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_710
timestamp 1626908933
transform 1 0 26900 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_142
timestamp 1626908933
transform 1 0 26688 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_864
timestamp 1626908933
transform 1 0 26688 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1063
timestamp 1626908933
transform 1 0 27552 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_462
timestamp 1626908933
transform 1 0 27552 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_568
timestamp 1626908933
transform 1 0 27456 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_211
timestamp 1626908933
transform 1 0 27456 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_871
timestamp 1626908933
transform 1 0 28272 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2838
timestamp 1626908933
transform 1 0 28272 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_867
timestamp 1626908933
transform 1 0 28944 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2834
timestamp 1626908933
transform 1 0 28944 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1449
timestamp 1626908933
transform 1 0 28080 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3416
timestamp 1626908933
transform 1 0 28080 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1533
timestamp 1626908933
transform 1 0 28848 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3468
timestamp 1626908933
transform 1 0 28848 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1677
timestamp 1626908933
transform 1 0 27888 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3644
timestamp 1626908933
transform 1 0 27888 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1448
timestamp 1626908933
transform 1 0 28080 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3415
timestamp 1626908933
transform 1 0 28080 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1650
timestamp 1626908933
transform 1 0 28272 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3617
timestamp 1626908933
transform 1 0 28272 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_85
timestamp 1626908933
transform 1 0 28560 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2052
timestamp 1626908933
transform 1 0 28560 0 1 12765
box -32 -32 32 32
use L1M1_PR  L1M1_PR_914
timestamp 1626908933
transform 1 0 29232 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_918
timestamp 1626908933
transform 1 0 29040 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2849
timestamp 1626908933
transform 1 0 29232 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2853
timestamp 1626908933
transform 1 0 29040 0 1 12321
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_38
timestamp 1626908933
transform 1 0 29300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_686
timestamp 1626908933
transform 1 0 29300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_38
timestamp 1626908933
transform 1 0 29300 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_686
timestamp 1626908933
transform 1 0 29300 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_196
timestamp 1626908933
transform 1 0 30048 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_797
timestamp 1626908933
transform 1 0 30048 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_382
timestamp 1626908933
transform 1 0 30240 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1373
timestamp 1626908933
transform 1 0 30240 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_95
timestamp 1626908933
transform 1 0 30000 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2030
timestamp 1626908933
transform 1 0 30000 0 1 12765
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_50
timestamp 1626908933
transform 1 0 30336 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_772
timestamp 1626908933
transform 1 0 30336 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_40
timestamp 1626908933
transform 1 0 27744 0 -1 13320
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_16
timestamp 1626908933
transform 1 0 27744 0 -1 13320
box -38 -49 2342 715
use M1M2_PR  M1M2_PR_3762
timestamp 1626908933
transform 1 0 30960 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1795
timestamp 1626908933
transform 1 0 30960 0 1 12839
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_606
timestamp 1626908933
transform 1 0 31104 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_8
timestamp 1626908933
transform 1 0 31104 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_381
timestamp 1626908933
transform 1 0 31488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1372
timestamp 1626908933
transform 1 0 31488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_210
timestamp 1626908933
transform 1 0 31680 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_567
timestamp 1626908933
transform 1 0 31680 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_816
timestamp 1626908933
transform 1 0 31584 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1807
timestamp 1626908933
transform 1 0 31584 0 -1 13320
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_14
timestamp 1626908933
transform 1 0 31700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_662
timestamp 1626908933
transform 1 0 31700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_14
timestamp 1626908933
transform 1 0 31700 0 1 12654
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_662
timestamp 1626908933
transform 1 0 31700 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_463
timestamp 1626908933
transform 1 0 31776 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1064
timestamp 1626908933
transform 1 0 31776 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3760
timestamp 1626908933
transform 1 0 32016 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1793
timestamp 1626908933
transform 1 0 32016 0 1 12839
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1808
timestamp 1626908933
transform 1 0 31968 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_817
timestamp 1626908933
transform 1 0 31968 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_209
timestamp 1626908933
transform 1 0 288 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_566
timestamp 1626908933
transform 1 0 288 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_464
timestamp 1626908933
transform 1 0 0 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1065
timestamp 1626908933
transform 1 0 0 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_818
timestamp 1626908933
transform 1 0 192 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_819
timestamp 1626908933
transform 1 0 384 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1809
timestamp 1626908933
transform 1 0 192 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1810
timestamp 1626908933
transform 1 0 384 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_9
timestamp 1626908933
transform 1 0 720 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1976
timestamp 1626908933
transform 1 0 720 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_11
timestamp 1626908933
transform 1 0 720 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1946
timestamp 1626908933
transform 1 0 720 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_5
timestamp 1626908933
transform -1 0 1344 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_13
timestamp 1626908933
transform -1 0 1344 0 1 13320
box -38 -49 902 715
use L1M1_PR  L1M1_PR_3807
timestamp 1626908933
transform 1 0 1104 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1872
timestamp 1626908933
transform 1 0 1104 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1943
timestamp 1626908933
transform 1 0 1200 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_8
timestamp 1626908933
transform 1 0 1200 0 1 13727
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1973
timestamp 1626908933
transform 1 0 1200 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_6
timestamp 1626908933
transform 1 0 1200 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3872
timestamp 1626908933
transform 1 0 1392 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1905
timestamp 1626908933
transform 1 0 1392 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1811
timestamp 1626908933
transform 1 0 1344 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_820
timestamp 1626908933
transform 1 0 1344 0 1 13320
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1286
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_638
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1286
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_638
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1940
timestamp 1626908933
transform 1 0 1584 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_5
timestamp 1626908933
transform 1 0 1584 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1971
timestamp 1626908933
transform 1 0 1488 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_4
timestamp 1626908933
transform 1 0 1488 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3804
timestamp 1626908933
transform 1 0 1872 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1869
timestamp 1626908933
transform 1 0 1872 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_1
timestamp 1626908933
transform -1 0 2304 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_9
timestamp 1626908933
transform -1 0 2304 0 1 13320
box -38 -49 902 715
use M1M2_PR  M1M2_PR_3300
timestamp 1626908933
transform 1 0 2640 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1333
timestamp 1626908933
transform 1 0 2640 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1371
timestamp 1626908933
transform 1 0 2304 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_380
timestamp 1626908933
transform 1 0 2304 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1148
timestamp 1626908933
transform 1 0 2400 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_550
timestamp 1626908933
transform 1 0 2400 0 1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1476
timestamp 1626908933
transform 1 0 3216 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3411
timestamp 1626908933
transform 1 0 3216 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1412
timestamp 1626908933
transform 1 0 2832 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3347
timestamp 1626908933
transform 1 0 2832 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1789
timestamp 1626908933
transform 1 0 3024 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3724
timestamp 1626908933
transform 1 0 3024 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1916
timestamp 1626908933
transform 1 0 3216 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3883
timestamp 1626908933
transform 1 0 3216 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1884
timestamp 1626908933
transform 1 0 3312 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3819
timestamp 1626908933
transform 1 0 3312 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1788
timestamp 1626908933
transform 1 0 3408 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3723
timestamp 1626908933
transform 1 0 3408 0 1 13727
box -29 -23 29 23
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_9
timestamp 1626908933
transform 1 0 2784 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_4
timestamp 1626908933
transform 1 0 2784 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_123
timestamp 1626908933
transform 1 0 3264 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_61
timestamp 1626908933
transform 1 0 3264 0 1 13320
box -38 -49 326 715
use M1M2_PR  M1M2_PR_3359
timestamp 1626908933
transform 1 0 3696 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1392
timestamp 1626908933
transform 1 0 3696 0 1 13431
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1262
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_614
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1262
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_614
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3629
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1694
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3565
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1598
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_630
timestamp 1626908933
transform 1 0 3552 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1352
timestamp 1626908933
transform 1 0 3552 0 1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3815
timestamp 1626908933
transform 1 0 4560 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3386
timestamp 1626908933
transform 1 0 4368 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1880
timestamp 1626908933
transform 1 0 4560 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1451
timestamp 1626908933
transform 1 0 4368 0 1 13579
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3879
timestamp 1626908933
transform 1 0 4560 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3335
timestamp 1626908933
transform 1 0 4272 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1912
timestamp 1626908933
transform 1 0 4560 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1368
timestamp 1626908933
transform 1 0 4272 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_47
timestamp 1626908933
transform 1 0 4320 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_22
timestamp 1626908933
transform 1 0 4320 0 1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3867
timestamp 1626908933
transform 1 0 4848 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3355
timestamp 1626908933
transform 1 0 4848 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1932
timestamp 1626908933
transform 1 0 4848 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1420
timestamp 1626908933
transform 1 0 4848 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1066
timestamp 1626908933
transform 1 0 4800 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_465
timestamp 1626908933
transform 1 0 4800 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_565
timestamp 1626908933
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_208
timestamp 1626908933
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1102
timestamp 1626908933
transform 1 0 5088 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_504
timestamp 1626908933
transform 1 0 5088 0 1 13320
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1363
timestamp 1626908933
transform 1 0 5520 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3330
timestamp 1626908933
transform 1 0 5520 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1446
timestamp 1626908933
transform 1 0 5520 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3381
timestamp 1626908933
transform 1 0 5520 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_9
timestamp 1626908933
transform 1 0 5472 0 1 13320
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_4
timestamp 1626908933
transform 1 0 5472 0 1 13320
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_432
timestamp 1626908933
transform 1 0 5808 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2399
timestamp 1626908933
transform 1 0 5808 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_428
timestamp 1626908933
transform 1 0 5712 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2363
timestamp 1626908933
transform 1 0 5712 0 1 13061
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_590
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1238
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_590
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1238
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1419
timestamp 1626908933
transform 1 0 5904 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3354
timestamp 1626908933
transform 1 0 5904 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_466
timestamp 1626908933
transform 1 0 7392 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1067
timestamp 1626908933
transform 1 0 7392 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_821
timestamp 1626908933
transform 1 0 7584 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1812
timestamp 1626908933
transform 1 0 7584 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1675
timestamp 1626908933
transform 1 0 7920 0 1 13505
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1676
timestamp 1626908933
transform 1 0 7920 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3642
timestamp 1626908933
transform 1 0 7920 0 1 13505
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3643
timestamp 1626908933
transform 1 0 7920 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1598
timestamp 1626908933
transform 1 0 7728 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1758
timestamp 1626908933
transform 1 0 7920 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3533
timestamp 1626908933
transform 1 0 7728 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3693
timestamp 1626908933
transform 1 0 7920 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1757
timestamp 1626908933
transform 1 0 8016 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3692
timestamp 1626908933
transform 1 0 8016 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_35
timestamp 1626908933
transform 1 0 7680 0 1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_10
timestamp 1626908933
transform 1 0 7680 0 1 13320
box -38 -49 2246 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1214
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_566
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1214
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_566
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3704
timestamp 1626908933
transform 1 0 8304 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1737
timestamp 1626908933
transform 1 0 8304 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3483
timestamp 1626908933
transform 1 0 9936 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1548
timestamp 1626908933
transform 1 0 9936 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3478
timestamp 1626908933
transform 1 0 9648 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1511
timestamp 1626908933
transform 1 0 9648 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1813
timestamp 1626908933
transform 1 0 9888 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_822
timestamp 1626908933
transform 1 0 9888 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_207
timestamp 1626908933
transform 1 0 9984 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_564
timestamp 1626908933
transform 1 0 9984 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_823
timestamp 1626908933
transform 1 0 10080 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1814
timestamp 1626908933
transform 1 0 10080 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_146
timestamp 1626908933
transform 1 0 10416 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2113
timestamp 1626908933
transform 1 0 10416 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_163
timestamp 1626908933
transform 1 0 10416 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1752
timestamp 1626908933
transform 1 0 10320 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2098
timestamp 1626908933
transform 1 0 10416 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3687
timestamp 1626908933
transform 1 0 10320 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_102
timestamp 1626908933
transform 1 0 10176 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_33
timestamp 1626908933
transform 1 0 10176 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_467
timestamp 1626908933
transform 1 0 10656 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1068
timestamp 1626908933
transform 1 0 10656 0 1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1462
timestamp 1626908933
transform 1 0 10704 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1463
timestamp 1626908933
transform 1 0 10704 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3429
timestamp 1626908933
transform 1 0 10704 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3430
timestamp 1626908933
transform 1 0 10704 0 1 13061
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_824
timestamp 1626908933
transform 1 0 10848 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1815
timestamp 1626908933
transform 1 0 10848 0 1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_890
timestamp 1626908933
transform 1 0 10992 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2825
timestamp 1626908933
transform 1 0 10992 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_18
timestamp 1626908933
transform -1 0 11328 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_80
timestamp 1626908933
transform -1 0 11328 0 1 13320
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1190
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_542
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1190
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_542
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2750
timestamp 1626908933
transform 1 0 11472 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_783
timestamp 1626908933
transform 1 0 11472 0 1 13209
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3482
timestamp 1626908933
transform 1 0 11088 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1547
timestamp 1626908933
transform 1 0 11088 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2749
timestamp 1626908933
transform 1 0 11184 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_814
timestamp 1626908933
transform 1 0 11184 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2749
timestamp 1626908933
transform 1 0 11472 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_782
timestamp 1626908933
transform 1 0 11472 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_17
timestamp 1626908933
transform 1 0 11904 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_78
timestamp 1626908933
transform 1 0 11904 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_468
timestamp 1626908933
transform 1 0 11712 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1069
timestamp 1626908933
transform 1 0 11712 0 1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_846
timestamp 1626908933
transform 1 0 11568 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2813
timestamp 1626908933
transform 1 0 11568 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_30
timestamp 1626908933
transform 1 0 11328 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_82
timestamp 1626908933
transform 1 0 11328 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_195
timestamp 1626908933
transform 1 0 12192 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_796
timestamp 1626908933
transform 1 0 12192 0 1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_61
timestamp 1626908933
transform 1 0 12240 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2028
timestamp 1626908933
transform 1 0 12240 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_68
timestamp 1626908933
transform 1 0 12144 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_888
timestamp 1626908933
transform 1 0 11952 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2003
timestamp 1626908933
transform 1 0 12144 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2823
timestamp 1626908933
transform 1 0 11952 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_471
timestamp 1626908933
transform 1 0 12384 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1193
timestamp 1626908933
transform 1 0 12384 0 1 13320
box -38 -49 806 715
use M1M2_PR  M1M2_PR_781
timestamp 1626908933
transform 1 0 13008 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2748
timestamp 1626908933
transform 1 0 13008 0 1 13209
box -32 -32 32 32
use L1M1_PR  L1M1_PR_64
timestamp 1626908933
transform 1 0 12912 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_813
timestamp 1626908933
transform 1 0 12912 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1999
timestamp 1626908933
transform 1 0 12912 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2748
timestamp 1626908933
transform 1 0 12912 0 1 13209
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_379
timestamp 1626908933
transform 1 0 13536 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1370
timestamp 1626908933
transform 1 0 13536 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_352
timestamp 1626908933
transform 1 0 13152 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_950
timestamp 1626908933
transform 1 0 13152 0 1 13320
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1166
timestamp 1626908933
transform 1 0 13700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_518
timestamp 1626908933
transform 1 0 13700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1166
timestamp 1626908933
transform 1 0 13700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_518
timestamp 1626908933
transform 1 0 13700 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1164
timestamp 1626908933
transform 1 0 13632 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_442
timestamp 1626908933
transform 1 0 13632 0 1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2746
timestamp 1626908933
transform 1 0 13872 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_811
timestamp 1626908933
transform 1 0 13872 0 1 13209
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2809
timestamp 1626908933
transform 1 0 14544 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_842
timestamp 1626908933
transform 1 0 14544 0 1 13209
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_795
timestamp 1626908933
transform 1 0 14400 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_194
timestamp 1626908933
transform 1 0 14400 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_931
timestamp 1626908933
transform 1 0 14592 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_333
timestamp 1626908933
transform 1 0 14592 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_206
timestamp 1626908933
transform 1 0 14976 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_563
timestamp 1626908933
transform 1 0 14976 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_193
timestamp 1626908933
transform 1 0 15072 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_794
timestamp 1626908933
transform 1 0 15072 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_378
timestamp 1626908933
transform 1 0 15264 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1369
timestamp 1626908933
transform 1 0 15264 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_840
timestamp 1626908933
transform 1 0 15312 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2807
timestamp 1626908933
transform 1 0 15312 0 1 13209
box -32 -32 32 32
use L1M1_PR  L1M1_PR_881
timestamp 1626908933
transform 1 0 15408 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_883
timestamp 1626908933
transform 1 0 15120 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2816
timestamp 1626908933
transform 1 0 15408 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2818
timestamp 1626908933
transform 1 0 15120 0 1 13209
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_409
timestamp 1626908933
transform 1 0 15360 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1131
timestamp 1626908933
transform 1 0 15360 0 1 13320
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_494
timestamp 1626908933
transform 1 0 16100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1142
timestamp 1626908933
transform 1 0 16100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_494
timestamp 1626908933
transform 1 0 16100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1142
timestamp 1626908933
transform 1 0 16100 0 1 13320
box -100 -49 100 49
use M1M2_PR  M1M2_PR_156
timestamp 1626908933
transform 1 0 15888 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_745
timestamp 1626908933
transform 1 0 16272 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2123
timestamp 1626908933
transform 1 0 15888 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2712
timestamp 1626908933
transform 1 0 16272 0 1 13431
box -32 -32 32 32
use L1M1_PR  L1M1_PR_171
timestamp 1626908933
transform 1 0 16176 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2106
timestamp 1626908933
transform 1 0 16176 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_2
timestamp 1626908933
transform 1 0 16128 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_8
timestamp 1626908933
transform 1 0 16128 0 1 13320
box -38 -49 518 715
use M1M2_PR  M1M2_PR_832
timestamp 1626908933
transform 1 0 16464 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2799
timestamp 1626908933
transform 1 0 16464 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_873
timestamp 1626908933
transform 1 0 16464 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_877
timestamp 1626908933
transform 1 0 16560 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2808
timestamp 1626908933
transform 1 0 16464 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2812
timestamp 1626908933
transform 1 0 16560 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_770
timestamp 1626908933
transform 1 0 16560 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2705
timestamp 1626908933
transform 1 0 16560 0 1 13431
box -29 -23 29 23
use M1M2_PR  M1M2_PR_749
timestamp 1626908933
transform 1 0 16464 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2716
timestamp 1626908933
transform 1 0 16464 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_658
timestamp 1626908933
transform 1 0 16560 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_775
timestamp 1626908933
transform 1 0 16368 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2593
timestamp 1626908933
transform 1 0 16560 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2710
timestamp 1626908933
transform 1 0 16368 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2814
timestamp 1626908933
transform 1 0 16848 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_879
timestamp 1626908933
transform 1 0 16848 0 1 13209
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_793
timestamp 1626908933
transform 1 0 16608 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_192
timestamp 1626908933
transform 1 0 16608 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1103
timestamp 1626908933
transform 1 0 16800 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_381
timestamp 1626908933
transform 1 0 16800 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_2
timestamp 1626908933
transform 1 0 17856 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_63
timestamp 1626908933
transform 1 0 17856 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_191
timestamp 1626908933
transform 1 0 17568 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_792
timestamp 1626908933
transform 1 0 17568 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_825
timestamp 1626908933
transform 1 0 17760 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1816
timestamp 1626908933
transform 1 0 17760 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2613
timestamp 1626908933
transform 1 0 17904 0 1 13135
box -32 -32 32 32
use M1M2_PR  M1M2_PR_646
timestamp 1626908933
transform 1 0 17904 0 1 13135
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2595
timestamp 1626908933
transform 1 0 18096 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_660
timestamp 1626908933
transform 1 0 18096 0 1 13431
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2612
timestamp 1626908933
transform 1 0 17904 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_645
timestamp 1626908933
transform 1 0 17904 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2007
timestamp 1626908933
transform 1 0 18096 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_72
timestamp 1626908933
transform 1 0 18096 0 1 13579
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2032
timestamp 1626908933
transform 1 0 18096 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_65
timestamp 1626908933
transform 1 0 18096 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_356
timestamp 1626908933
transform 1 0 18144 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1078
timestamp 1626908933
transform 1 0 18144 0 1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2592
timestamp 1626908933
transform 1 0 18384 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_657
timestamp 1626908933
transform 1 0 18384 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2596
timestamp 1626908933
transform 1 0 18576 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2588
timestamp 1626908933
transform 1 0 18672 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_661
timestamp 1626908933
transform 1 0 18576 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_653
timestamp 1626908933
transform 1 0 18672 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2616
timestamp 1626908933
transform 1 0 18480 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_649
timestamp 1626908933
transform 1 0 18480 0 1 13061
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1118
timestamp 1626908933
transform 1 0 18500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_470
timestamp 1626908933
transform 1 0 18500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1118
timestamp 1626908933
transform 1 0 18500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_470
timestamp 1626908933
transform 1 0 18500 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2594
timestamp 1626908933
transform 1 0 18960 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2591
timestamp 1626908933
transform 1 0 18768 0 1 13135
box -29 -23 29 23
use L1M1_PR  L1M1_PR_659
timestamp 1626908933
transform 1 0 18960 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_656
timestamp 1626908933
transform 1 0 18768 0 1 13135
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2615
timestamp 1626908933
transform 1 0 18864 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_648
timestamp 1626908933
transform 1 0 18864 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2718
timestamp 1626908933
transform 1 0 19056 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2651
timestamp 1626908933
transform 1 0 19056 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2614
timestamp 1626908933
transform 1 0 18864 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_751
timestamp 1626908933
transform 1 0 19056 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_684
timestamp 1626908933
transform 1 0 19056 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_647
timestamp 1626908933
transform 1 0 18864 0 1 13431
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1070
timestamp 1626908933
transform 1 0 18912 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_469
timestamp 1626908933
transform 1 0 18912 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_10
timestamp 1626908933
transform -1 0 19488 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_72
timestamp 1626908933
transform -1 0 19488 0 1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2712
timestamp 1626908933
transform 1 0 19152 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2590
timestamp 1626908933
transform 1 0 19152 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2024
timestamp 1626908933
transform 1 0 19344 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_777
timestamp 1626908933
transform 1 0 19152 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_655
timestamp 1626908933
transform 1 0 19152 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_89
timestamp 1626908933
transform 1 0 19344 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2046
timestamp 1626908933
transform 1 0 19344 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_79
timestamp 1626908933
transform 1 0 19344 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2635
timestamp 1626908933
transform 1 0 19536 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_700
timestamp 1626908933
transform 1 0 19536 0 1 13431
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2045
timestamp 1626908933
transform 1 0 19440 0 1 13135
box -32 -32 32 32
use M1M2_PR  M1M2_PR_78
timestamp 1626908933
transform 1 0 19440 0 1 13135
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1817
timestamp 1626908933
transform 1 0 19872 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_826
timestamp 1626908933
transform 1 0 19872 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_83
timestamp 1626908933
transform 1 0 19488 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_31
timestamp 1626908933
transform 1 0 19488 0 1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2022
timestamp 1626908933
transform 1 0 20112 0 1 13135
box -29 -23 29 23
use L1M1_PR  L1M1_PR_87
timestamp 1626908933
transform 1 0 20112 0 1 13135
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2823
timestamp 1626908933
transform 1 0 20112 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2042
timestamp 1626908933
transform 1 0 19920 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_856
timestamp 1626908933
transform 1 0 20112 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_75
timestamp 1626908933
transform 1 0 19920 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1071
timestamp 1626908933
transform 1 0 20064 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_470
timestamp 1626908933
transform 1 0 20064 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_562
timestamp 1626908933
transform 1 0 19968 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_205
timestamp 1626908933
transform 1 0 19968 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_827
timestamp 1626908933
transform 1 0 20256 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1818
timestamp 1626908933
transform 1 0 20256 0 1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_81
timestamp 1626908933
transform 1 0 20400 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2016
timestamp 1626908933
transform 1 0 20400 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_92
timestamp 1626908933
transform 1 0 20352 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_23
timestamp 1626908933
transform 1 0 20352 0 1 13320
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1094
timestamp 1626908933
transform 1 0 20900 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_446
timestamp 1626908933
transform 1 0 20900 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1094
timestamp 1626908933
transform 1 0 20900 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_446
timestamp 1626908933
transform 1 0 20900 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_801
timestamp 1626908933
transform 1 0 20832 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_203
timestamp 1626908933
transform 1 0 20832 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_82
timestamp 1626908933
transform -1 0 21504 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_20
timestamp 1626908933
transform -1 0 21504 0 1 13320
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2834
timestamp 1626908933
transform 1 0 21264 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_899
timestamp 1626908933
transform 1 0 21264 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3419
timestamp 1626908933
transform 1 0 21360 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1452
timestamp 1626908933
transform 1 0 21360 0 1 13061
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1072
timestamp 1626908933
transform 1 0 21504 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_471
timestamp 1626908933
transform 1 0 21504 0 1 13320
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3675
timestamp 1626908933
transform 1 0 21936 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1740
timestamp 1626908933
transform 1 0 21936 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2650
timestamp 1626908933
transform 1 0 21744 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_683
timestamp 1626908933
transform 1 0 21744 0 1 13431
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1819
timestamp 1626908933
transform 1 0 21696 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_828
timestamp 1626908933
transform 1 0 21696 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_36
timestamp 1626908933
transform -1 0 22272 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_105
timestamp 1626908933
transform -1 0 22272 0 1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3472
timestamp 1626908933
transform 1 0 22320 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1537
timestamp 1626908933
transform 1 0 22320 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2503
timestamp 1626908933
transform 1 0 22128 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2119
timestamp 1626908933
transform 1 0 22224 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_568
timestamp 1626908933
transform 1 0 22128 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_184
timestamp 1626908933
transform 1 0 22224 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2135
timestamp 1626908933
transform 1 0 22320 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_168
timestamp 1626908933
transform 1 0 22320 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_791
timestamp 1626908933
transform 1 0 22272 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_190
timestamp 1626908933
transform 1 0 22272 0 1 13320
box -38 -49 230 715
use L1M1_PR  L1M1_PR_567
timestamp 1626908933
transform 1 0 22896 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2502
timestamp 1626908933
transform 1 0 22896 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_31
timestamp 1626908933
transform 1 0 22848 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_93
timestamp 1626908933
transform 1 0 22848 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_176
timestamp 1626908933
transform 1 0 22464 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_774
timestamp 1626908933
transform 1 0 22464 0 1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2951
timestamp 1626908933
transform 1 0 23088 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1016
timestamp 1626908933
transform 1 0 23088 0 1 13727
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2531
timestamp 1626908933
transform 1 0 22992 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_564
timestamp 1626908933
transform 1 0 22992 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1368
timestamp 1626908933
transform 1 0 23136 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_377
timestamp 1626908933
transform 1 0 23136 0 1 13320
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1070
timestamp 1626908933
transform 1 0 23300 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_422
timestamp 1626908933
transform 1 0 23300 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1070
timestamp 1626908933
transform 1 0 23300 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_422
timestamp 1626908933
transform 1 0 23300 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3674
timestamp 1626908933
transform 1 0 23280 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1739
timestamp 1626908933
transform 1 0 23280 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_953
timestamp 1626908933
transform 1 0 23760 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2920
timestamp 1626908933
transform 1 0 23760 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_233
timestamp 1626908933
transform 1 0 23232 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_955
timestamp 1626908933
transform 1 0 23232 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_189
timestamp 1626908933
transform 1 0 24000 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_790
timestamp 1626908933
transform 1 0 24000 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_376
timestamp 1626908933
transform 1 0 24192 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1367
timestamp 1626908933
transform 1 0 24192 0 1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2955
timestamp 1626908933
transform 1 0 24432 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2949
timestamp 1626908933
transform 1 0 24240 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2122
timestamp 1626908933
transform 1 0 24528 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1020
timestamp 1626908933
transform 1 0 24432 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1014
timestamp 1626908933
transform 1 0 24240 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_187
timestamp 1626908933
transform 1 0 24528 0 1 13579
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2139
timestamp 1626908933
transform 1 0 24336 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_172
timestamp 1626908933
transform 1 0 24336 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_87
timestamp 1626908933
transform 1 0 24288 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_26
timestamp 1626908933
transform 1 0 24288 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_134
timestamp 1626908933
transform 1 0 24576 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_732
timestamp 1626908933
transform 1 0 24576 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_204
timestamp 1626908933
transform 1 0 24960 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_561
timestamp 1626908933
transform 1 0 24960 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_123
timestamp 1626908933
transform 1 0 25152 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_721
timestamp 1626908933
transform 1 0 25152 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_375
timestamp 1626908933
transform 1 0 25056 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1366
timestamp 1626908933
transform 1 0 25056 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2922
timestamp 1626908933
transform 1 0 25488 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_955
timestamp 1626908933
transform 1 0 25488 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1365
timestamp 1626908933
transform 1 0 25536 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_374
timestamp 1626908933
transform 1 0 25536 0 1 13320
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1046
timestamp 1626908933
transform 1 0 25700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_398
timestamp 1626908933
transform 1 0 25700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1046
timestamp 1626908933
transform 1 0 25700 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_398
timestamp 1626908933
transform 1 0 25700 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2953
timestamp 1626908933
transform 1 0 25776 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1018
timestamp 1626908933
transform 1 0 25776 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1820
timestamp 1626908933
transform 1 0 25632 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_829
timestamp 1626908933
transform 1 0 25632 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_92
timestamp 1626908933
transform -1 0 26016 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_30
timestamp 1626908933
transform -1 0 26016 0 1 13320
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2957
timestamp 1626908933
transform 1 0 25872 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2688
timestamp 1626908933
transform 1 0 25968 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1022
timestamp 1626908933
transform 1 0 25872 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_753
timestamp 1626908933
transform 1 0 25968 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3461
timestamp 1626908933
transform 1 0 25872 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1494
timestamp 1626908933
transform 1 0 25872 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1364
timestamp 1626908933
transform 1 0 26016 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_373
timestamp 1626908933
transform 1 0 26016 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2924
timestamp 1626908933
transform 1 0 26256 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2694
timestamp 1626908933
transform 1 0 26064 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_957
timestamp 1626908933
transform 1 0 26256 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_727
timestamp 1626908933
transform 1 0 26064 0 1 13653
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_704
timestamp 1626908933
transform 1 0 26112 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_106
timestamp 1626908933
transform 1 0 26112 0 1 13320
box -38 -49 422 715
use M1M2_PR  M1M2_PR_175
timestamp 1626908933
transform 1 0 26640 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1686
timestamp 1626908933
transform 1 0 26544 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2142
timestamp 1626908933
transform 1 0 26640 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3653
timestamp 1626908933
transform 1 0 26544 0 1 13727
box -32 -32 32 32
use L1M1_PR  L1M1_PR_191
timestamp 1626908933
transform 1 0 26640 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2126
timestamp 1626908933
transform 1 0 26640 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_372
timestamp 1626908933
transform 1 0 27264 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1363
timestamp 1626908933
transform 1 0 27264 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1651
timestamp 1626908933
transform 1 0 27504 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3618
timestamp 1626908933
transform 1 0 27504 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1581
timestamp 1626908933
transform 1 0 27408 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3516
timestamp 1626908933
transform 1 0 27408 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_158
timestamp 1626908933
transform 1 0 26496 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_880
timestamp 1626908933
transform 1 0 26496 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_43
timestamp 1626908933
transform 1 0 27360 0 1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_18
timestamp 1626908933
transform 1 0 27360 0 1 13320
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_1534
timestamp 1626908933
transform 1 0 27792 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3469
timestamp 1626908933
transform 1 0 27792 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1732
timestamp 1626908933
transform 1 0 28176 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3667
timestamp 1626908933
transform 1 0 28176 0 1 12987
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_374
timestamp 1626908933
transform 1 0 28100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1022
timestamp 1626908933
transform 1 0 28100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_374
timestamp 1626908933
transform 1 0 28100 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1022
timestamp 1626908933
transform 1 0 28100 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1734
timestamp 1626908933
transform 1 0 27696 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3669
timestamp 1626908933
transform 1 0 27696 0 1 13579
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1649
timestamp 1626908933
transform 1 0 28272 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3616
timestamp 1626908933
transform 1 0 28272 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2125
timestamp 1626908933
transform 1 0 29520 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_190
timestamp 1626908933
transform 1 0 29520 0 1 13431
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_789
timestamp 1626908933
transform 1 0 30048 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_188
timestamp 1626908933
transform 1 0 30048 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_641
timestamp 1626908933
transform 1 0 29568 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_43
timestamp 1626908933
transform 1 0 29568 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_560
timestamp 1626908933
transform 1 0 29952 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_203
timestamp 1626908933
transform 1 0 29952 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1362
timestamp 1626908933
transform 1 0 30240 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_371
timestamp 1626908933
transform 1 0 30240 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_771
timestamp 1626908933
transform 1 0 30336 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_49
timestamp 1626908933
transform 1 0 30336 0 1 13320
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_998
timestamp 1626908933
transform 1 0 30500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_350
timestamp 1626908933
transform 1 0 30500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_998
timestamp 1626908933
transform 1 0 30500 0 1 13320
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_350
timestamp 1626908933
transform 1 0 30500 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1361
timestamp 1626908933
transform 1 0 31104 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_370
timestamp 1626908933
transform 1 0 31104 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_735
timestamp 1626908933
transform 1 0 31200 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_13
timestamp 1626908933
transform 1 0 31200 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1821
timestamp 1626908933
transform 1 0 31968 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_830
timestamp 1626908933
transform 1 0 31968 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_187
timestamp 1626908933
transform 1 0 0 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_788
timestamp 1626908933
transform 1 0 0 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1877
timestamp 1626908933
transform 1 0 48 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3844
timestamp 1626908933
transform 1 0 48 0 1 14245
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_325
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_973
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_325
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_973
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_713
timestamp 1626908933
transform 1 0 192 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1435
timestamp 1626908933
transform 1 0 192 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1360
timestamp 1626908933
transform 1 0 960 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_369
timestamp 1626908933
transform 1 0 960 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1173
timestamp 1626908933
transform 1 0 1056 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_575
timestamp 1626908933
transform 1 0 1056 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1401
timestamp 1626908933
transform 1 0 1440 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_679
timestamp 1626908933
transform 1 0 1440 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_368
timestamp 1626908933
transform 1 0 2208 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1359
timestamp 1626908933
transform 1 0 2208 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3
timestamp 1626908933
transform 1 0 2160 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1970
timestamp 1626908933
transform 1 0 2160 0 1 13875
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3
timestamp 1626908933
transform 1 0 2160 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1938
timestamp 1626908933
transform 1 0 2160 0 1 13875
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_202
timestamp 1626908933
transform 1 0 2496 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_559
timestamp 1626908933
transform 1 0 2496 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_472
timestamp 1626908933
transform 1 0 2304 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1073
timestamp 1626908933
transform 1 0 2304 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1358
timestamp 1626908933
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_367
timestamp 1626908933
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1376
timestamp 1626908933
transform 1 0 2688 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_654
timestamp 1626908933
transform 1 0 2688 0 -1 14652
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_949
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_301
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_949
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_301
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1135
timestamp 1626908933
transform 1 0 3456 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_537
timestamp 1626908933
transform 1 0 3456 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3334
timestamp 1626908933
transform 1 0 4272 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1367
timestamp 1626908933
transform 1 0 4272 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_787
timestamp 1626908933
transform 1 0 3840 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_186
timestamp 1626908933
transform 1 0 3840 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1351
timestamp 1626908933
transform 1 0 4032 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_629
timestamp 1626908933
transform 1 0 4032 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_366
timestamp 1626908933
transform 1 0 4800 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1357
timestamp 1626908933
transform 1 0 4800 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1911
timestamp 1626908933
transform 1 0 4560 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3878
timestamp 1626908933
transform 1 0 4560 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1812
timestamp 1626908933
transform 1 0 5136 0 1 14467
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3779
timestamp 1626908933
transform 1 0 5136 0 1 14467
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_277
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_925
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_277
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_925
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_510
timestamp 1626908933
transform 1 0 4896 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1108
timestamp 1626908933
transform 1 0 4896 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_21
timestamp 1626908933
transform 1 0 5280 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_46
timestamp 1626908933
transform 1 0 5280 0 -1 14652
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1362
timestamp 1626908933
transform 1 0 5520 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1910
timestamp 1626908933
transform 1 0 5424 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3329
timestamp 1626908933
transform 1 0 5520 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3877
timestamp 1626908933
transform 1 0 5424 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1909
timestamp 1626908933
transform 1 0 5424 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3876
timestamp 1626908933
transform 1 0 5424 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1449
timestamp 1626908933
transform 1 0 5328 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1877
timestamp 1626908933
transform 1 0 5520 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3384
timestamp 1626908933
transform 1 0 5328 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3812
timestamp 1626908933
transform 1 0 5520 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3738
timestamp 1626908933
transform 1 0 6000 0 1 14467
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1803
timestamp 1626908933
transform 1 0 6000 0 1 14467
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1822
timestamp 1626908933
transform 1 0 5952 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_831
timestamp 1626908933
transform 1 0 5952 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1074
timestamp 1626908933
transform 1 0 5760 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_473
timestamp 1626908933
transform 1 0 5760 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_62
timestamp 1626908933
transform 1 0 6048 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_131
timestamp 1626908933
transform 1 0 6048 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_30
timestamp 1626908933
transform -1 0 7104 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_5
timestamp 1626908933
transform -1 0 7104 0 -1 14652
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3380
timestamp 1626908933
transform 1 0 6192 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1445
timestamp 1626908933
transform 1 0 6192 0 1 14097
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3842
timestamp 1626908933
transform 1 0 6288 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1875
timestamp 1626908933
transform 1 0 6288 0 1 14245
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1823
timestamp 1626908933
transform 1 0 6528 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_832
timestamp 1626908933
transform 1 0 6528 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1365
timestamp 1626908933
transform 1 0 6864 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3332
timestamp 1626908933
transform 1 0 6864 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1448
timestamp 1626908933
transform 1 0 6864 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3383
timestamp 1626908933
transform 1 0 6864 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3388
timestamp 1626908933
transform 1 0 7056 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1453
timestamp 1626908933
transform 1 0 7056 0 1 13875
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3337
timestamp 1626908933
transform 1 0 7056 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1370
timestamp 1626908933
transform 1 0 7056 0 1 13875
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3387
timestamp 1626908933
transform 1 0 7056 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1452
timestamp 1626908933
transform 1 0 7056 0 1 14393
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3336
timestamp 1626908933
transform 1 0 7056 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1369
timestamp 1626908933
transform 1 0 7056 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1824
timestamp 1626908933
transform 1 0 7104 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_833
timestamp 1626908933
transform 1 0 7104 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_35
timestamp 1626908933
transform -1 0 7488 0 -1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_96
timestamp 1626908933
transform -1 0 7488 0 -1 14652
box -38 -49 326 715
use M1M2_PR  M1M2_PR_900
timestamp 1626908933
transform 1 0 7248 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1946
timestamp 1626908933
transform 1 0 7248 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2867
timestamp 1626908933
transform 1 0 7248 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3913
timestamp 1626908933
transform 1 0 7248 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_947
timestamp 1626908933
transform 1 0 7344 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1721
timestamp 1626908933
transform 1 0 7440 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2882
timestamp 1626908933
transform 1 0 7344 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3656
timestamp 1626908933
transform 1 0 7440 0 1 14393
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_201
timestamp 1626908933
transform 1 0 7488 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_558
timestamp 1626908933
transform 1 0 7488 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1637
timestamp 1626908933
transform 1 0 7536 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3604
timestamp 1626908933
transform 1 0 7536 0 1 14393
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_253
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_901
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_253
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_901
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_469
timestamp 1626908933
transform 1 0 7584 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1067
timestamp 1626908933
transform 1 0 7584 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_804
timestamp 1626908933
transform 1 0 8112 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2771
timestamp 1626908933
transform 1 0 8112 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1674
timestamp 1626908933
transform 1 0 7920 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3641
timestamp 1626908933
transform 1 0 7920 0 1 14245
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1755
timestamp 1626908933
transform 1 0 8208 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1909
timestamp 1626908933
transform 1 0 8112 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3690
timestamp 1626908933
transform 1 0 8208 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3844
timestamp 1626908933
transform 1 0 8112 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_1
timestamp 1626908933
transform -1 0 8352 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_0
timestamp 1626908933
transform -1 0 8352 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_474
timestamp 1626908933
transform 1 0 8352 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1075
timestamp 1626908933
transform 1 0 8352 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_834
timestamp 1626908933
transform 1 0 8544 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1825
timestamp 1626908933
transform 1 0 8544 0 -1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1714
timestamp 1626908933
transform 1 0 8592 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3649
timestamp 1626908933
transform 1 0 8592 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_516
timestamp 1626908933
transform 1 0 8880 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_838
timestamp 1626908933
transform 1 0 8880 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2451
timestamp 1626908933
transform 1 0 8880 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2773
timestamp 1626908933
transform 1 0 8880 0 1 14097
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_441
timestamp 1626908933
transform 1 0 9120 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1039
timestamp 1626908933
transform 1 0 9120 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_0
timestamp 1626908933
transform 1 0 8640 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2b_1  sky130_fd_sc_hs__nand2b_1_5
timestamp 1626908933
transform 1 0 8640 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_835
timestamp 1626908933
transform 1 0 9504 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1826
timestamp 1626908933
transform 1 0 9504 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1510
timestamp 1626908933
transform 1 0 9648 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3477
timestamp 1626908933
transform 1 0 9648 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_676
timestamp 1626908933
transform 1 0 9840 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_989
timestamp 1626908933
transform 1 0 9936 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1597
timestamp 1626908933
transform 1 0 9648 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2611
timestamp 1626908933
transform 1 0 9840 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2924
timestamp 1626908933
transform 1 0 9936 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3532
timestamp 1626908933
transform 1 0 9648 0 1 14097
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_516
timestamp 1626908933
transform 1 0 9984 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1238
timestamp 1626908933
transform 1 0 9984 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_30
timestamp 1626908933
transform -1 0 9984 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_92
timestamp 1626908933
transform -1 0 9984 0 -1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2610
timestamp 1626908933
transform 1 0 10320 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_675
timestamp 1626908933
transform 1 0 10320 0 1 13875
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2627
timestamp 1626908933
transform 1 0 10320 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_660
timestamp 1626908933
transform 1 0 10320 0 1 13875
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_877
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_229
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_877
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_229
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2626
timestamp 1626908933
transform 1 0 10320 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_659
timestamp 1626908933
transform 1 0 10320 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_932
timestamp 1626908933
transform 1 0 10608 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2899
timestamp 1626908933
transform 1 0 10608 0 1 14245
box -32 -32 32 32
use L1M1_PR  L1M1_PR_674
timestamp 1626908933
transform 1 0 10800 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2609
timestamp 1626908933
transform 1 0 10800 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_34
timestamp 1626908933
transform 1 0 10752 0 -1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_96
timestamp 1626908933
transform 1 0 10752 0 -1 14652
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2922
timestamp 1626908933
transform 1 0 10992 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_987
timestamp 1626908933
transform 1 0 10992 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_84
timestamp 1626908933
transform 1 0 11040 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_32
timestamp 1626908933
transform 1 0 11040 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_475
timestamp 1626908933
transform 1 0 11424 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1076
timestamp 1626908933
transform 1 0 11424 0 -1 14652
box -38 -49 230 715
use L1M1_PR  L1M1_PR_886
timestamp 1626908933
transform 1 0 11376 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2821
timestamp 1626908933
transform 1 0 11376 0 1 13875
box -29 -23 29 23
use M1M2_PR  M1M2_PR_845
timestamp 1626908933
transform 1 0 11568 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2812
timestamp 1626908933
transform 1 0 11568 0 1 14245
box -32 -32 32 32
use L1M1_PR  L1M1_PR_71
timestamp 1626908933
transform 1 0 11568 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_889
timestamp 1626908933
transform 1 0 11760 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2006
timestamp 1626908933
transform 1 0 11568 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2824
timestamp 1626908933
transform 1 0 11760 0 1 14245
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_5
timestamp 1626908933
transform -1 0 12192 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_44
timestamp 1626908933
transform -1 0 12192 0 -1 14652
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2828
timestamp 1626908933
transform 1 0 12048 0 1 13801
box -29 -23 29 23
use L1M1_PR  L1M1_PR_893
timestamp 1626908933
transform 1 0 12048 0 1 13801
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2818
timestamp 1626908933
transform 1 0 12048 0 1 13801
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2027
timestamp 1626908933
transform 1 0 12240 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_851
timestamp 1626908933
transform 1 0 12048 0 1 13801
box -32 -32 32 32
use M1M2_PR  M1M2_PR_60
timestamp 1626908933
transform 1 0 12240 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2829
timestamp 1626908933
transform 1 0 11952 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_894
timestamp 1626908933
transform 1 0 11952 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2817
timestamp 1626908933
transform 1 0 12048 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_850
timestamp 1626908933
transform 1 0 12048 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1077
timestamp 1626908933
transform 1 0 12192 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_476
timestamp 1626908933
transform 1 0 12192 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_200
timestamp 1626908933
transform 1 0 12480 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_557
timestamp 1626908933
transform 1 0 12480 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_836
timestamp 1626908933
transform 1 0 12384 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1827
timestamp 1626908933
transform 1 0 12384 0 -1 14652
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_205
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_853
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_205
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_853
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_364
timestamp 1626908933
transform 1 0 12576 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_962
timestamp 1626908933
transform 1 0 12576 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_780
timestamp 1626908933
transform 1 0 13008 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2747
timestamp 1626908933
transform 1 0 13008 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_812
timestamp 1626908933
transform 1 0 13008 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_887
timestamp 1626908933
transform 1 0 13104 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2747
timestamp 1626908933
transform 1 0 13008 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2822
timestamp 1626908933
transform 1 0 13104 0 1 14245
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_22
timestamp 1626908933
transform 1 0 12960 0 -1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_84
timestamp 1626908933
transform 1 0 12960 0 -1 14652
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2820
timestamp 1626908933
transform 1 0 13200 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_885
timestamp 1626908933
transform 1 0 13200 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2811
timestamp 1626908933
transform 1 0 13200 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2810
timestamp 1626908933
transform 1 0 13200 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_844
timestamp 1626908933
transform 1 0 13200 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_843
timestamp 1626908933
transform 1 0 13200 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1356
timestamp 1626908933
transform 1 0 13440 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_365
timestamp 1626908933
transform 1 0 13440 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_786
timestamp 1626908933
transform 1 0 13248 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_185
timestamp 1626908933
transform 1 0 13248 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_441
timestamp 1626908933
transform 1 0 13536 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1163
timestamp 1626908933
transform 1 0 13536 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_43
timestamp 1626908933
transform 1 0 14304 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_4
timestamp 1626908933
transform 1 0 14304 0 -1 14652
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2819
timestamp 1626908933
transform 1 0 14544 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_884
timestamp 1626908933
transform 1 0 14544 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2808
timestamp 1626908933
transform 1 0 14544 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2019
timestamp 1626908933
transform 1 0 14160 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_841
timestamp 1626908933
transform 1 0 14544 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_52
timestamp 1626908933
transform 1 0 14160 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_839
timestamp 1626908933
transform 1 0 15312 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2806
timestamp 1626908933
transform 1 0 15312 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_882
timestamp 1626908933
transform 1 0 14736 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2817
timestamp 1626908933
transform 1 0 14736 0 1 14097
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_181
timestamp 1626908933
transform 1 0 14900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_829
timestamp 1626908933
transform 1 0 14900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_181
timestamp 1626908933
transform 1 0 14900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_829
timestamp 1626908933
transform 1 0 14900 0 1 13986
box -100 -49 100 49
use L1M1_PR  L1M1_PR_59
timestamp 1626908933
transform 1 0 14832 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1994
timestamp 1626908933
transform 1 0 14832 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_422
timestamp 1626908933
transform 1 0 14880 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1144
timestamp 1626908933
transform 1 0 14880 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_364
timestamp 1626908933
transform 1 0 15648 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1355
timestamp 1626908933
transform 1 0 15648 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_656
timestamp 1626908933
transform 1 0 15696 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2623
timestamp 1626908933
transform 1 0 15696 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_363
timestamp 1626908933
transform 1 0 16128 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1354
timestamp 1626908933
transform 1 0 16128 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_68
timestamp 1626908933
transform 1 0 16272 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2035
timestamp 1626908933
transform 1 0 16272 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_392
timestamp 1626908933
transform 1 0 16224 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1114
timestamp 1626908933
transform 1 0 16224 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_305
timestamp 1626908933
transform 1 0 15744 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_903
timestamp 1626908933
transform 1 0 15744 0 -1 14652
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_805
timestamp 1626908933
transform 1 0 17300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_157
timestamp 1626908933
transform 1 0 17300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_805
timestamp 1626908933
transform 1 0 17300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_157
timestamp 1626908933
transform 1 0 17300 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1353
timestamp 1626908933
transform 1 0 16992 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_362
timestamp 1626908933
transform 1 0 16992 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_878
timestamp 1626908933
transform 1 0 17088 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_280
timestamp 1626908933
transform 1 0 17088 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2816
timestamp 1626908933
transform 1 0 17520 0 1 13801
box -32 -32 32 32
use M1M2_PR  M1M2_PR_849
timestamp 1626908933
transform 1 0 17520 0 1 13801
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_556
timestamp 1626908933
transform 1 0 17472 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_199
timestamp 1626908933
transform 1 0 17472 0 -1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2008
timestamp 1626908933
transform 1 0 17616 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_73
timestamp 1626908933
transform 1 0 17616 0 1 14393
box -29 -23 29 23
use M1M2_PR  M1M2_PR_653
timestamp 1626908933
transform 1 0 17808 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2620
timestamp 1626908933
transform 1 0 17808 0 1 13875
box -32 -32 32 32
use L1M1_PR  L1M1_PR_665
timestamp 1626908933
transform 1 0 17808 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2600
timestamp 1626908933
transform 1 0 17808 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_662
timestamp 1626908933
transform 1 0 17808 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2597
timestamp 1626908933
transform 1 0 17808 0 1 14097
box -29 -23 29 23
use M1M2_PR  M1M2_PR_652
timestamp 1626908933
transform 1 0 17808 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2619
timestamp 1626908933
transform 1 0 17808 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_664
timestamp 1626908933
transform 1 0 17808 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2599
timestamp 1626908933
transform 1 0 17808 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_64
timestamp 1626908933
transform 1 0 18096 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2031
timestamp 1626908933
transform 1 0 18096 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_80
timestamp 1626908933
transform 1 0 18192 0 1 14171
box -29 -23 29 23
use L1M1_PR  L1M1_PR_785
timestamp 1626908933
transform 1 0 17904 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2015
timestamp 1626908933
transform 1 0 18192 0 1 14171
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2720
timestamp 1626908933
transform 1 0 17904 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_13
timestamp 1626908933
transform 1 0 18144 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_36
timestamp 1626908933
transform 1 0 18144 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_4
timestamp 1626908933
transform 1 0 17568 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_10
timestamp 1626908933
transform 1 0 17568 0 -1 14652
box -38 -49 614 715
use M1M2_PR  M1M2_PR_651
timestamp 1626908933
transform 1 0 18288 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2618
timestamp 1626908933
transform 1 0 18288 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_72
timestamp 1626908933
transform 1 0 18672 0 1 14171
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2039
timestamp 1626908933
transform 1 0 18672 0 1 14171
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_477
timestamp 1626908933
transform 1 0 18912 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1078
timestamp 1626908933
transform 1 0 18912 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_750
timestamp 1626908933
transform 1 0 19056 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2717
timestamp 1626908933
transform 1 0 19056 0 1 14097
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_837
timestamp 1626908933
transform 1 0 19104 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1828
timestamp 1626908933
transform 1 0 19104 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_28
timestamp 1626908933
transform -1 0 19872 0 -1 14652
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_13
timestamp 1626908933
transform -1 0 19872 0 -1 14652
box -38 -49 710 715
use L1M1_PR  L1M1_PR_2711
timestamp 1626908933
transform 1 0 19248 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_776
timestamp 1626908933
transform 1 0 19248 0 1 14097
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2722
timestamp 1626908933
transform 1 0 19344 0 1 14467
box -32 -32 32 32
use M1M2_PR  M1M2_PR_755
timestamp 1626908933
transform 1 0 19344 0 1 14467
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_781
timestamp 1626908933
transform 1 0 19700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_133
timestamp 1626908933
transform 1 0 19700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_781
timestamp 1626908933
transform 1 0 19700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_133
timestamp 1626908933
transform 1 0 19700 0 1 13986
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2718
timestamp 1626908933
transform 1 0 19536 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2716
timestamp 1626908933
transform 1 0 19440 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_783
timestamp 1626908933
transform 1 0 19536 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_781
timestamp 1626908933
transform 1 0 19440 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2012
timestamp 1626908933
transform 1 0 19728 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_77
timestamp 1626908933
transform 1 0 19728 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_184
timestamp 1626908933
transform 1 0 19872 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_785
timestamp 1626908933
transform 1 0 19872 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_855
timestamp 1626908933
transform 1 0 20112 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2822
timestamp 1626908933
transform 1 0 20112 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_308
timestamp 1626908933
transform 1 0 20064 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1030
timestamp 1626908933
transform 1 0 20064 0 -1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_860
timestamp 1626908933
transform 1 0 20976 0 1 13801
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2827
timestamp 1626908933
transform 1 0 20976 0 1 13801
box -32 -32 32 32
use L1M1_PR  L1M1_PR_905
timestamp 1626908933
transform 1 0 20688 0 1 13801
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2840
timestamp 1626908933
transform 1 0 20688 0 1 13801
box -29 -23 29 23
use M1M2_PR  M1M2_PR_859
timestamp 1626908933
transform 1 0 20976 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2826
timestamp 1626908933
transform 1 0 20976 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_900
timestamp 1626908933
transform 1 0 20880 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_904
timestamp 1626908933
transform 1 0 20976 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2835
timestamp 1626908933
transform 1 0 20880 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2839
timestamp 1626908933
transform 1 0 20976 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_20
timestamp 1626908933
transform 1 0 20832 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_82
timestamp 1626908933
transform 1 0 20832 0 -1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2843
timestamp 1626908933
transform 1 0 21168 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_908
timestamp 1626908933
transform 1 0 21168 0 1 14393
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1352
timestamp 1626908933
transform 1 0 21216 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_361
timestamp 1626908933
transform 1 0 21216 0 -1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2841
timestamp 1626908933
transform 1 0 21264 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_906
timestamp 1626908933
transform 1 0 21264 0 1 13875
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2829
timestamp 1626908933
transform 1 0 21264 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2828
timestamp 1626908933
transform 1 0 21264 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2132
timestamp 1626908933
transform 1 0 21360 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_862
timestamp 1626908933
transform 1 0 21264 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_861
timestamp 1626908933
transform 1 0 21264 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_165
timestamp 1626908933
transform 1 0 21360 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2838
timestamp 1626908933
transform 1 0 21552 0 1 13801
box -29 -23 29 23
use L1M1_PR  L1M1_PR_903
timestamp 1626908933
transform 1 0 21552 0 1 13801
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2916
timestamp 1626908933
transform 1 0 21840 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_949
timestamp 1626908933
transform 1 0 21840 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2649
timestamp 1626908933
transform 1 0 21744 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_682
timestamp 1626908933
transform 1 0 21744 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2634
timestamp 1626908933
transform 1 0 21840 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_699
timestamp 1626908933
transform 1 0 21840 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2114
timestamp 1626908933
transform 1 0 21744 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_179
timestamp 1626908933
transform 1 0 21744 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2915
timestamp 1626908933
transform 1 0 21840 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_948
timestamp 1626908933
transform 1 0 21840 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_77
timestamp 1626908933
transform 1 0 21696 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_8
timestamp 1626908933
transform 1 0 21696 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_195
timestamp 1626908933
transform 1 0 21312 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_793
timestamp 1626908933
transform 1 0 21312 0 -1 14652
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_757
timestamp 1626908933
transform 1 0 22100 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_109
timestamp 1626908933
transform 1 0 22100 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_757
timestamp 1626908933
transform 1 0 22100 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_109
timestamp 1626908933
transform 1 0 22100 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_198
timestamp 1626908933
transform 1 0 22464 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_555
timestamp 1626908933
transform 1 0 22464 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_478
timestamp 1626908933
transform 1 0 22176 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1079
timestamp 1626908933
transform 1 0 22176 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_838
timestamp 1626908933
transform 1 0 22368 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1829
timestamp 1626908933
transform 1 0 22368 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_183
timestamp 1626908933
transform 1 0 22560 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_784
timestamp 1626908933
transform 1 0 22560 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_360
timestamp 1626908933
transform 1 0 22752 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1351
timestamp 1626908933
transform 1 0 22752 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_174
timestamp 1626908933
transform 1 0 22848 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_772
timestamp 1626908933
transform 1 0 22848 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_563
timestamp 1626908933
transform 1 0 22992 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2530
timestamp 1626908933
transform 1 0 22992 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_566
timestamp 1626908933
transform 1 0 23376 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1009
timestamp 1626908933
transform 1 0 23280 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1010
timestamp 1626908933
transform 1 0 23184 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2501
timestamp 1626908933
transform 1 0 23376 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2944
timestamp 1626908933
transform 1 0 23280 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2945
timestamp 1626908933
transform 1 0 23184 0 1 13875
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_182
timestamp 1626908933
transform 1 0 23616 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_783
timestamp 1626908933
transform 1 0 23616 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_359
timestamp 1626908933
transform 1 0 23808 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1350
timestamp 1626908933
transform 1 0 23808 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_952
timestamp 1626908933
transform 1 0 23760 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2919
timestamp 1626908933
transform 1 0 23760 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1015
timestamp 1626908933
transform 1 0 23568 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2950
timestamp 1626908933
transform 1 0 23568 0 1 14393
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_33
timestamp 1626908933
transform 1 0 23232 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_95
timestamp 1626908933
transform 1 0 23232 0 -1 14652
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_733
timestamp 1626908933
transform 1 0 24500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_85
timestamp 1626908933
transform 1 0 24500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_733
timestamp 1626908933
transform 1 0 24500 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_85
timestamp 1626908933
transform 1 0 24500 0 1 13986
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2138
timestamp 1626908933
transform 1 0 24336 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_171
timestamp 1626908933
transform 1 0 24336 0 1 14097
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_942
timestamp 1626908933
transform 1 0 23904 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_220
timestamp 1626908933
transform 1 0 23904 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1349
timestamp 1626908933
transform 1 0 24672 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_358
timestamp 1626908933
transform 1 0 24672 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_909
timestamp 1626908933
transform 1 0 24768 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_187
timestamp 1626908933
transform 1 0 24768 0 -1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_954
timestamp 1626908933
transform 1 0 25488 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2921
timestamp 1626908933
transform 1 0 25488 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_20
timestamp 1626908933
transform 1 0 25536 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_59
timestamp 1626908933
transform 1 0 25536 0 -1 14652
box -38 -49 614 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_6
timestamp 1626908933
transform 1 0 26112 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_58
timestamp 1626908933
transform 1 0 26112 0 -1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_186
timestamp 1626908933
transform 1 0 26160 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1013
timestamp 1626908933
transform 1 0 25968 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1017
timestamp 1626908933
transform 1 0 25776 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2121
timestamp 1626908933
transform 1 0 26160 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2948
timestamp 1626908933
transform 1 0 25968 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2952
timestamp 1626908933
transform 1 0 25776 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1798
timestamp 1626908933
transform 1 0 26736 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3765
timestamp 1626908933
transform 1 0 26736 0 1 13875
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_61
timestamp 1626908933
transform 1 0 26900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_709
timestamp 1626908933
transform 1 0 26900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_61
timestamp 1626908933
transform 1 0 26900 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_709
timestamp 1626908933
transform 1 0 26900 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_197
timestamp 1626908933
transform 1 0 27456 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_554
timestamp 1626908933
transform 1 0 27456 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_479
timestamp 1626908933
transform 1 0 27264 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1080
timestamp 1626908933
transform 1 0 27264 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_170
timestamp 1626908933
transform 1 0 27408 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2137
timestamp 1626908933
transform 1 0 27408 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1486
timestamp 1626908933
transform 1 0 27600 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3421
timestamp 1626908933
transform 1 0 27600 0 1 14393
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_157
timestamp 1626908933
transform 1 0 26496 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_879
timestamp 1626908933
transform 1 0 26496 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_58
timestamp 1626908933
transform 1 0 27552 0 -1 14652
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_12
timestamp 1626908933
transform 1 0 27552 0 -1 14652
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3389
timestamp 1626908933
transform 1 0 27984 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1454
timestamp 1626908933
transform 1 0 27984 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3370
timestamp 1626908933
transform 1 0 28464 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3338
timestamp 1626908933
transform 1 0 27696 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2344
timestamp 1626908933
transform 1 0 27888 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1403
timestamp 1626908933
transform 1 0 28464 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1371
timestamp 1626908933
transform 1 0 27696 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_377
timestamp 1626908933
transform 1 0 27888 0 1 14245
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_685
timestamp 1626908933
transform 1 0 29300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_37
timestamp 1626908933
transform 1 0 29300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_685
timestamp 1626908933
transform 1 0 29300 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_37
timestamp 1626908933
transform 1 0 29300 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1348
timestamp 1626908933
transform 1 0 30240 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_357
timestamp 1626908933
transform 1 0 30240 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_770
timestamp 1626908933
transform 1 0 30336 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_48
timestamp 1626908933
transform 1 0 30336 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_605
timestamp 1626908933
transform 1 0 31104 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_7
timestamp 1626908933
transform 1 0 31104 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_356
timestamp 1626908933
transform 1 0 31488 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1347
timestamp 1626908933
transform 1 0 31488 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_196
timestamp 1626908933
transform 1 0 31680 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_553
timestamp 1626908933
transform 1 0 31680 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_839
timestamp 1626908933
transform 1 0 31584 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1830
timestamp 1626908933
transform 1 0 31584 0 -1 14652
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_13
timestamp 1626908933
transform 1 0 31700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_661
timestamp 1626908933
transform 1 0 31700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_13
timestamp 1626908933
transform 1 0 31700 0 1 13986
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_661
timestamp 1626908933
transform 1 0 31700 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_480
timestamp 1626908933
transform 1 0 31776 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1081
timestamp 1626908933
transform 1 0 31776 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3763
timestamp 1626908933
transform 1 0 32016 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1796
timestamp 1626908933
transform 1 0 32016 0 1 13875
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1831
timestamp 1626908933
transform 1 0 31968 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_840
timestamp 1626908933
transform 1 0 31968 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3780
timestamp 1626908933
transform 1 0 48 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1813
timestamp 1626908933
transform 1 0 48 0 1 15059
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1832
timestamp 1626908933
transform 1 0 192 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_841
timestamp 1626908933
transform 1 0 192 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1833
timestamp 1626908933
transform 1 0 384 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_842
timestamp 1626908933
transform 1 0 384 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_552
timestamp 1626908933
transform 1 0 288 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_195
timestamp 1626908933
transform 1 0 288 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1082
timestamp 1626908933
transform 1 0 0 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_481
timestamp 1626908933
transform 1 0 0 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_8
timestamp 1626908933
transform 1 0 720 0 1 15133
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1975
timestamp 1626908933
transform 1 0 720 0 1 15133
box -32 -32 32 32
use L1M1_PR  L1M1_PR_10
timestamp 1626908933
transform 1 0 720 0 1 15133
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1874
timestamp 1626908933
transform 1 0 720 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1945
timestamp 1626908933
transform 1 0 720 0 1 15133
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3809
timestamp 1626908933
transform 1 0 720 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_6
timestamp 1626908933
transform 1 0 480 0 1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_14
timestamp 1626908933
transform 1 0 480 0 1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_482
timestamp 1626908933
transform 1 0 1344 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1083
timestamp 1626908933
transform 1 0 1344 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1904
timestamp 1626908933
transform 1 0 1392 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3871
timestamp 1626908933
transform 1 0 1392 0 1 14911
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1808
timestamp 1626908933
transform 1 0 1008 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3743
timestamp 1626908933
transform 1 0 1008 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1807
timestamp 1626908933
transform 1 0 1680 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1871
timestamp 1626908933
transform 1 0 1680 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3742
timestamp 1626908933
transform 1 0 1680 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3806
timestamp 1626908933
transform 1 0 1680 0 1 14985
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_637
timestamp 1626908933
transform 1 0 1700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1285
timestamp 1626908933
transform 1 0 1700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_637
timestamp 1626908933
transform 1 0 1700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1285
timestamp 1626908933
transform 1 0 1700 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_0
timestamp 1626908933
transform 1 0 1536 0 1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_8
timestamp 1626908933
transform 1 0 1536 0 1 14652
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1937
timestamp 1626908933
transform 1 0 2160 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2
timestamp 1626908933
transform 1 0 2160 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3299
timestamp 1626908933
transform 1 0 2640 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1969
timestamp 1626908933
transform 1 0 2160 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1332
timestamp 1626908933
transform 1 0 2640 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2
timestamp 1626908933
transform 1 0 2160 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1147
timestamp 1626908933
transform 1 0 2400 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_549
timestamp 1626908933
transform 1 0 2400 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_483
timestamp 1626908933
transform 1 0 2784 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1084
timestamp 1626908933
transform 1 0 2784 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1337
timestamp 1626908933
transform 1 0 3120 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3304
timestamp 1626908933
transform 1 0 3120 0 1 15207
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1416
timestamp 1626908933
transform 1 0 3024 0 1 15207
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3351
timestamp 1626908933
transform 1 0 3024 0 1 15207
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1915
timestamp 1626908933
transform 1 0 3216 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3882
timestamp 1626908933
transform 1 0 3216 0 1 14911
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1411
timestamp 1626908933
transform 1 0 3408 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1885
timestamp 1626908933
transform 1 0 3216 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3346
timestamp 1626908933
transform 1 0 3408 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3820
timestamp 1626908933
transform 1 0 3216 0 1 14911
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_536
timestamp 1626908933
transform 1 0 3456 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1134
timestamp 1626908933
transform 1 0 3456 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_20
timestamp 1626908933
transform -1 0 3456 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_45
timestamp 1626908933
transform -1 0 3456 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_484
timestamp 1626908933
transform 1 0 3840 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1085
timestamp 1626908933
transform 1 0 3840 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_843
timestamp 1626908933
transform 1 0 4032 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1834
timestamp 1626908933
transform 1 0 4032 0 1 14652
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1261
timestamp 1626908933
transform 1 0 4100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_613
timestamp 1626908933
transform 1 0 4100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1261
timestamp 1626908933
transform 1 0 4100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_613
timestamp 1626908933
transform 1 0 4100 0 1 14652
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3741
timestamp 1626908933
transform 1 0 4080 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1806
timestamp 1626908933
transform 1 0 4080 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2454
timestamp 1626908933
transform 1 0 4368 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_519
timestamp 1626908933
transform 1 0 4368 0 1 14911
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3333
timestamp 1626908933
transform 1 0 4272 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1366
timestamp 1626908933
transform 1 0 4272 0 1 14837
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_0
timestamp 1626908933
transform 1 0 4128 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_25
timestamp 1626908933
transform 1 0 4128 0 1 14652
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1450
timestamp 1626908933
transform 1 0 4464 0 1 14837
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3385
timestamp 1626908933
transform 1 0 4464 0 1 14837
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_194
timestamp 1626908933
transform 1 0 4992 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_551
timestamp 1626908933
transform 1 0 4992 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_181
timestamp 1626908933
transform 1 0 5088 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_782
timestamp 1626908933
transform 1 0 5088 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_604
timestamp 1626908933
transform 1 0 5280 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1326
timestamp 1626908933
transform 1 0 5280 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_518
timestamp 1626908933
transform 1 0 4608 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1116
timestamp 1626908933
transform 1 0 4608 0 1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_521
timestamp 1626908933
transform 1 0 6096 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1339
timestamp 1626908933
transform 1 0 5616 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2488
timestamp 1626908933
transform 1 0 6096 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3306
timestamp 1626908933
transform 1 0 5616 0 1 14541
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1417
timestamp 1626908933
transform 1 0 5616 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3352
timestamp 1626908933
transform 1 0 5616 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_520
timestamp 1626908933
transform 1 0 6096 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2487
timestamp 1626908933
transform 1 0 6096 0 1 14911
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_492
timestamp 1626908933
transform 1 0 6048 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1090
timestamp 1626908933
transform 1 0 6048 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_355
timestamp 1626908933
transform 1 0 6432 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1346
timestamp 1626908933
transform 1 0 6432 0 1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_518
timestamp 1626908933
transform 1 0 6768 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2453
timestamp 1626908933
transform 1 0 6768 0 1 14541
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_589
timestamp 1626908933
transform 1 0 6500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1237
timestamp 1626908933
transform 1 0 6500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_589
timestamp 1626908933
transform 1 0 6500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1237
timestamp 1626908933
transform 1 0 6500 0 1 14652
box -100 -49 100 49
use L1M1_PR  L1M1_PR_517
timestamp 1626908933
transform 1 0 7152 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2452
timestamp 1626908933
transform 1 0 7152 0 1 14541
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_576
timestamp 1626908933
transform 1 0 6528 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1298
timestamp 1626908933
transform 1 0 6528 0 1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3640
timestamp 1626908933
transform 1 0 7920 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1673
timestamp 1626908933
transform 1 0 7920 0 1 14911
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_781
timestamp 1626908933
transform 1 0 7296 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_180
timestamp 1626908933
transform 1 0 7296 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1066
timestamp 1626908933
transform 1 0 7488 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_468
timestamp 1626908933
transform 1 0 7488 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1278
timestamp 1626908933
transform 1 0 7872 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_556
timestamp 1626908933
transform 1 0 7872 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_354
timestamp 1626908933
transform 1 0 8640 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1345
timestamp 1626908933
transform 1 0 8640 0 1 14652
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_565
timestamp 1626908933
transform 1 0 8900 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1213
timestamp 1626908933
transform 1 0 8900 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_565
timestamp 1626908933
transform 1 0 8900 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1213
timestamp 1626908933
transform 1 0 8900 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_537
timestamp 1626908933
transform 1 0 9120 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1259
timestamp 1626908933
transform 1 0 9120 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_446
timestamp 1626908933
transform 1 0 8736 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1044
timestamp 1626908933
transform 1 0 8736 0 1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2928
timestamp 1626908933
transform 1 0 9552 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_993
timestamp 1626908933
transform 1 0 9552 0 1 14541
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1835
timestamp 1626908933
transform 1 0 9888 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_844
timestamp 1626908933
transform 1 0 9888 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_550
timestamp 1626908933
transform 1 0 9984 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_193
timestamp 1626908933
transform 1 0 9984 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1020
timestamp 1626908933
transform 1 0 10080 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_422
timestamp 1626908933
transform 1 0 10080 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1237
timestamp 1626908933
transform 1 0 10464 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_515
timestamp 1626908933
transform 1 0 10464 0 1 14652
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2927
timestamp 1626908933
transform 1 0 10896 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_992
timestamp 1626908933
transform 1 0 10896 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2903
timestamp 1626908933
transform 1 0 10992 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_936
timestamp 1626908933
transform 1 0 10992 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_395
timestamp 1626908933
transform 1 0 11328 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_993
timestamp 1626908933
transform 1 0 11328 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_353
timestamp 1626908933
transform 1 0 11232 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1344
timestamp 1626908933
transform 1 0 11232 0 1 14652
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_541
timestamp 1626908933
transform 1 0 11300 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1189
timestamp 1626908933
transform 1 0 11300 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_541
timestamp 1626908933
transform 1 0 11300 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1189
timestamp 1626908933
transform 1 0 11300 0 1 14652
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1461
timestamp 1626908933
transform 1 0 12144 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3428
timestamp 1626908933
transform 1 0 12144 0 1 14541
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1546
timestamp 1626908933
transform 1 0 12144 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3481
timestamp 1626908933
transform 1 0 12144 0 1 14541
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_485
timestamp 1626908933
transform 1 0 11712 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1207
timestamp 1626908933
transform 1 0 11712 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_352
timestamp 1626908933
transform 1 0 12480 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_845
timestamp 1626908933
transform 1 0 12576 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1343
timestamp 1626908933
transform 1 0 12480 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1836
timestamp 1626908933
transform 1 0 12576 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1464
timestamp 1626908933
transform 1 0 12720 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1465
timestamp 1626908933
transform 1 0 12720 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3431
timestamp 1626908933
transform 1 0 12720 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3432
timestamp 1626908933
transform 1 0 12720 0 1 14541
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1550
timestamp 1626908933
transform 1 0 12720 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3485
timestamp 1626908933
transform 1 0 12720 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1669
timestamp 1626908933
transform 1 0 13008 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3636
timestamp 1626908933
transform 1 0 13008 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1725
timestamp 1626908933
transform 1 0 13200 0 1 15133
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3692
timestamp 1626908933
transform 1 0 13200 0 1 15133
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1750
timestamp 1626908933
transform 1 0 13104 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3685
timestamp 1626908933
transform 1 0 13104 0 1 14985
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_517
timestamp 1626908933
transform 1 0 13700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1165
timestamp 1626908933
transform 1 0 13700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_517
timestamp 1626908933
transform 1 0 13700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1165
timestamp 1626908933
transform 1 0 13700 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_33
timestamp 1626908933
transform 1 0 12672 0 1 14652
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_9
timestamp 1626908933
transform 1 0 12672 0 1 14652
box -38 -49 2342 715
use L1M1_PR  L1M1_PR_3484
timestamp 1626908933
transform 1 0 14352 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1549
timestamp 1626908933
transform 1 0 14352 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2018
timestamp 1626908933
transform 1 0 14160 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_51
timestamp 1626908933
transform 1 0 14160 0 1 14763
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1993
timestamp 1626908933
transform 1 0 14928 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_58
timestamp 1626908933
transform 1 0 14928 0 1 14763
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1837
timestamp 1626908933
transform 1 0 15456 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_846
timestamp 1626908933
transform 1 0 15456 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_918
timestamp 1626908933
transform 1 0 15072 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_320
timestamp 1626908933
transform 1 0 15072 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_549
timestamp 1626908933
transform 1 0 14976 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_192
timestamp 1626908933
transform 1 0 14976 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_655
timestamp 1626908933
transform 1 0 15696 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2622
timestamp 1626908933
transform 1 0 15696 0 1 15207
box -32 -32 32 32
use L1M1_PR  L1M1_PR_667
timestamp 1626908933
transform 1 0 15696 0 1 15207
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2602
timestamp 1626908933
transform 1 0 15696 0 1 15207
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1141
timestamp 1626908933
transform 1 0 16100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_493
timestamp 1626908933
transform 1 0 16100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1141
timestamp 1626908933
transform 1 0 16100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_493
timestamp 1626908933
transform 1 0 16100 0 1 14652
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2107
timestamp 1626908933
transform 1 0 15888 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_172
timestamp 1626908933
transform 1 0 15888 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2122
timestamp 1626908933
transform 1 0 15888 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_155
timestamp 1626908933
transform 1 0 15888 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1086
timestamp 1626908933
transform 1 0 16032 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_485
timestamp 1626908933
transform 1 0 16032 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_103
timestamp 1626908933
transform -1 0 16032 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_34
timestamp 1626908933
transform -1 0 16032 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_847
timestamp 1626908933
transform 1 0 16224 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1838
timestamp 1626908933
transform 1 0 16224 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_67
timestamp 1626908933
transform 1 0 16272 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2034
timestamp 1626908933
transform 1 0 16272 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_748
timestamp 1626908933
transform 1 0 16464 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2715
timestamp 1626908933
transform 1 0 16464 0 1 14763
box -32 -32 32 32
use L1M1_PR  L1M1_PR_74
timestamp 1626908933
transform 1 0 16464 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_774
timestamp 1626908933
transform 1 0 16464 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2009
timestamp 1626908933
transform 1 0 16464 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2709
timestamp 1626908933
transform 1 0 16464 0 1 14763
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_91
timestamp 1626908933
transform -1 0 16800 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_22
timestamp 1626908933
transform -1 0 16800 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1102
timestamp 1626908933
transform 1 0 16800 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_380
timestamp 1626908933
transform 1 0 16800 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_351
timestamp 1626908933
transform 1 0 17568 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1342
timestamp 1626908933
transform 1 0 17568 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1901
timestamp 1626908933
transform 1 0 17712 0 1 15133
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3868
timestamp 1626908933
transform 1 0 17712 0 1 15133
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_350
timestamp 1626908933
transform 1 0 18048 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1341
timestamp 1626908933
transform 1 0 18048 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_355
timestamp 1626908933
transform 1 0 18144 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1077
timestamp 1626908933
transform 1 0 18144 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_268
timestamp 1626908933
transform 1 0 17664 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_866
timestamp 1626908933
transform 1 0 17664 0 1 14652
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_469
timestamp 1626908933
transform 1 0 18500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1117
timestamp 1626908933
transform 1 0 18500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_469
timestamp 1626908933
transform 1 0 18500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1117
timestamp 1626908933
transform 1 0 18500 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_179
timestamp 1626908933
transform 1 0 18912 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_780
timestamp 1626908933
transform 1 0 18912 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_757
timestamp 1626908933
transform 1 0 19056 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2724
timestamp 1626908933
transform 1 0 19056 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_349
timestamp 1626908933
transform 1 0 19104 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1340
timestamp 1626908933
transform 1 0 19104 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1049
timestamp 1626908933
transform 1 0 19200 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_327
timestamp 1626908933
transform 1 0 19200 0 1 14652
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2018
timestamp 1626908933
transform 1 0 19824 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_83
timestamp 1626908933
transform 1 0 19824 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2041
timestamp 1626908933
transform 1 0 19920 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_74
timestamp 1626908933
transform 1 0 19920 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1029
timestamp 1626908933
transform 1 0 20064 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_307
timestamp 1626908933
transform 1 0 20064 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_548
timestamp 1626908933
transform 1 0 19968 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_191
timestamp 1626908933
transform 1 0 19968 0 1 14652
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1093
timestamp 1626908933
transform 1 0 20900 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_445
timestamp 1626908933
transform 1 0 20900 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1093
timestamp 1626908933
transform 1 0 20900 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_445
timestamp 1626908933
transform 1 0 20900 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1339
timestamp 1626908933
transform 1 0 20832 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_348
timestamp 1626908933
transform 1 0 20832 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_800
timestamp 1626908933
transform 1 0 20928 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_202
timestamp 1626908933
transform 1 0 20928 0 1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3475
timestamp 1626908933
transform 1 0 21072 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1540
timestamp 1626908933
transform 1 0 21072 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3624
timestamp 1626908933
transform 1 0 21552 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1657
timestamp 1626908933
transform 1 0 21552 0 1 14911
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1005
timestamp 1626908933
transform 1 0 21312 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_283
timestamp 1626908933
transform 1 0 21312 0 1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3422
timestamp 1626908933
transform 1 0 21936 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1455
timestamp 1626908933
transform 1 0 21936 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_783
timestamp 1626908933
transform 1 0 22080 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_185
timestamp 1626908933
transform 1 0 22080 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_347
timestamp 1626908933
transform 1 0 22464 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1338
timestamp 1626908933
transform 1 0 22464 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_167
timestamp 1626908933
transform 1 0 22320 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2134
timestamp 1626908933
transform 1 0 22320 0 1 14763
box -32 -32 32 32
use L1M1_PR  L1M1_PR_182
timestamp 1626908933
transform 1 0 22608 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2117
timestamp 1626908933
transform 1 0 22608 0 1 14763
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1691
timestamp 1626908933
transform 1 0 22992 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3658
timestamp 1626908933
transform 1 0 22992 0 1 14985
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_421
timestamp 1626908933
transform 1 0 23300 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1069
timestamp 1626908933
transform 1 0 23300 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_421
timestamp 1626908933
transform 1 0 23300 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1069
timestamp 1626908933
transform 1 0 23300 0 1 14652
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1586
timestamp 1626908933
transform 1 0 23472 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3521
timestamp 1626908933
transform 1 0 23472 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1900
timestamp 1626908933
transform 1 0 23856 0 1 15133
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3867
timestamp 1626908933
transform 1 0 23856 0 1 15133
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1737
timestamp 1626908933
transform 1 0 24432 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3672
timestamp 1626908933
transform 1 0 24432 0 1 14911
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_486
timestamp 1626908933
transform 1 0 24768 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1087
timestamp 1626908933
transform 1 0 24768 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1498
timestamp 1626908933
transform 1 0 24624 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1499
timestamp 1626908933
transform 1 0 24624 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3465
timestamp 1626908933
transform 1 0 24624 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3466
timestamp 1626908933
transform 1 0 24624 0 1 14541
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1585
timestamp 1626908933
transform 1 0 24720 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3520
timestamp 1626908933
transform 1 0 24720 0 1 14911
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_41
timestamp 1626908933
transform -1 0 24768 0 1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_16
timestamp 1626908933
transform -1 0 24768 0 1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_190
timestamp 1626908933
transform 1 0 24960 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_547
timestamp 1626908933
transform 1 0 24960 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_487
timestamp 1626908933
transform 1 0 25056 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1088
timestamp 1626908933
transform 1 0 25056 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1496
timestamp 1626908933
transform 1 0 25392 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1497
timestamp 1626908933
transform 1 0 25392 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3463
timestamp 1626908933
transform 1 0 25392 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3464
timestamp 1626908933
transform 1 0 25392 0 1 14541
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1584
timestamp 1626908933
transform 1 0 25296 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3519
timestamp 1626908933
transform 1 0 25296 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1583
timestamp 1626908933
transform 1 0 25584 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1736
timestamp 1626908933
transform 1 0 25584 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3518
timestamp 1626908933
transform 1 0 25584 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3671
timestamp 1626908933
transform 1 0 25584 0 1 14911
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_397
timestamp 1626908933
transform 1 0 25700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1045
timestamp 1626908933
transform 1 0 25700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_397
timestamp 1626908933
transform 1 0 25700 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1045
timestamp 1626908933
transform 1 0 25700 0 1 14652
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1801
timestamp 1626908933
transform 1 0 25872 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3768
timestamp 1626908933
transform 1 0 25872 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1687
timestamp 1626908933
transform 1 0 26448 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3654
timestamp 1626908933
transform 1 0 26448 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1654
timestamp 1626908933
transform 1 0 27312 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3621
timestamp 1626908933
transform 1 0 27312 0 1 14837
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_178
timestamp 1626908933
transform 1 0 27456 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_779
timestamp 1626908933
transform 1 0 27456 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_169
timestamp 1626908933
transform 1 0 27408 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2136
timestamp 1626908933
transform 1 0 27408 0 1 14763
box -32 -32 32 32
use L1M1_PR  L1M1_PR_185
timestamp 1626908933
transform 1 0 27408 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2120
timestamp 1626908933
transform 1 0 27408 0 1 14763
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_346
timestamp 1626908933
transform 1 0 27648 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1337
timestamp 1626908933
transform 1 0 27648 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_42
timestamp 1626908933
transform 1 0 25248 0 1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_17
timestamp 1626908933
transform 1 0 25248 0 1 14652
box -38 -49 2246 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1021
timestamp 1626908933
transform 1 0 28100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_373
timestamp 1626908933
transform 1 0 28100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1021
timestamp 1626908933
transform 1 0 28100 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_373
timestamp 1626908933
transform 1 0 28100 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_848
timestamp 1626908933
transform 1 0 27744 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_126
timestamp 1626908933
transform 1 0 27744 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1336
timestamp 1626908933
transform 1 0 28896 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_345
timestamp 1626908933
transform 1 0 28896 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_660
timestamp 1626908933
transform 1 0 28512 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_62
timestamp 1626908933
transform 1 0 28512 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_814
timestamp 1626908933
transform 1 0 28992 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_92
timestamp 1626908933
transform 1 0 28992 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_488
timestamp 1626908933
transform 1 0 29760 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1089
timestamp 1626908933
transform 1 0 29760 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_189
timestamp 1626908933
transform 1 0 29952 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_546
timestamp 1626908933
transform 1 0 29952 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_177
timestamp 1626908933
transform 1 0 30048 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_778
timestamp 1626908933
transform 1 0 30048 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_360
timestamp 1626908933
transform 1 0 29904 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2327
timestamp 1626908933
transform 1 0 29904 0 1 14541
box -32 -32 32 32
use L1M1_PR  L1M1_PR_383
timestamp 1626908933
transform 1 0 29904 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2318
timestamp 1626908933
transform 1 0 29904 0 1 14541
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1335
timestamp 1626908933
transform 1 0 30240 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_344
timestamp 1626908933
transform 1 0 30240 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_769
timestamp 1626908933
transform 1 0 30336 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_47
timestamp 1626908933
transform 1 0 30336 0 1 14652
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_997
timestamp 1626908933
transform 1 0 30500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_349
timestamp 1626908933
transform 1 0 30500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_997
timestamp 1626908933
transform 1 0 30500 0 1 14652
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_349
timestamp 1626908933
transform 1 0 30500 0 1 14652
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1334
timestamp 1626908933
transform 1 0 31104 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_343
timestamp 1626908933
transform 1 0 31104 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_734
timestamp 1626908933
transform 1 0 31200 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_12
timestamp 1626908933
transform 1 0 31200 0 1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3766
timestamp 1626908933
transform 1 0 32016 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1799
timestamp 1626908933
transform 1 0 32016 0 1 15207
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1839
timestamp 1626908933
transform 1 0 31968 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_848
timestamp 1626908933
transform 1 0 31968 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1842
timestamp 1626908933
transform 1 0 192 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_851
timestamp 1626908933
transform 1 0 192 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1094
timestamp 1626908933
transform 1 0 0 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_777
timestamp 1626908933
transform 1 0 0 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_493
timestamp 1626908933
transform 1 0 0 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_176
timestamp 1626908933
transform 1 0 0 0 -1 15984
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_972
timestamp 1626908933
transform 1 0 500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_324
timestamp 1626908933
transform 1 0 500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_972
timestamp 1626908933
transform 1 0 500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_324
timestamp 1626908933
transform 1 0 500 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_538
timestamp 1626908933
transform 1 0 288 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_181
timestamp 1626908933
transform 1 0 288 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_574
timestamp 1626908933
transform 1 0 1056 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1172
timestamp 1626908933
transform 1 0 1056 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_342
timestamp 1626908933
transform 1 0 960 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1333
timestamp 1626908933
transform 1 0 960 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_712
timestamp 1626908933
transform 1 0 192 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1434
timestamp 1626908933
transform 1 0 192 0 -1 15984
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_636
timestamp 1626908933
transform 1 0 1700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1284
timestamp 1626908933
transform 1 0 1700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_636
timestamp 1626908933
transform 1 0 1700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1284
timestamp 1626908933
transform 1 0 1700 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1332
timestamp 1626908933
transform 1 0 2208 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_341
timestamp 1626908933
transform 1 0 2208 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1090
timestamp 1626908933
transform 1 0 2304 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_489
timestamp 1626908933
transform 1 0 2304 0 -1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3931
timestamp 1626908933
transform 1 0 2448 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1964
timestamp 1626908933
transform 1 0 2448 0 1 15725
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_545
timestamp 1626908933
transform 1 0 2496 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_188
timestamp 1626908933
transform 1 0 2496 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3869
timestamp 1626908933
transform 1 0 2640 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1934
timestamp 1626908933
transform 1 0 2640 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_678
timestamp 1626908933
transform 1 0 1440 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1400
timestamp 1626908933
transform 1 0 1440 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_46
timestamp 1626908933
transform -1 0 3072 0 1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_0
timestamp 1626908933
transform -1 0 3072 0 1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_7
timestamp 1626908933
transform 1 0 2592 0 -1 15984
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_2
timestamp 1626908933
transform 1 0 2592 0 -1 15984
box -38 -49 1958 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_300
timestamp 1626908933
transform 1 0 2900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_948
timestamp 1626908933
transform 1 0 2900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_300
timestamp 1626908933
transform 1 0 2900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_948
timestamp 1626908933
transform 1 0 2900 0 1 15318
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1415
timestamp 1626908933
transform 1 0 3024 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3350
timestamp 1626908933
transform 1 0 3024 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1336
timestamp 1626908933
transform 1 0 3120 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3303
timestamp 1626908933
transform 1 0 3120 0 1 15651
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_612
timestamp 1626908933
transform 1 0 4100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1260
timestamp 1626908933
transform 1 0 4100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_612
timestamp 1626908933
transform 1 0 4100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1260
timestamp 1626908933
transform 1 0 4100 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_517
timestamp 1626908933
transform 1 0 4608 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1115
timestamp 1626908933
transform 1 0 4608 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_340
timestamp 1626908933
transform 1 0 4512 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1331
timestamp 1626908933
transform 1 0 4512 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1805
timestamp 1626908933
transform 1 0 4368 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3740
timestamp 1626908933
transform 1 0 4368 0 1 15577
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_180
timestamp 1626908933
transform 1 0 4992 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_537
timestamp 1626908933
transform 1 0 4992 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_339
timestamp 1626908933
transform 1 0 4992 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1330
timestamp 1626908933
transform 1 0 4992 0 -1 15984
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_276
timestamp 1626908933
transform 1 0 5300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_924
timestamp 1626908933
transform 1 0 5300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_276
timestamp 1626908933
transform 1 0 5300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_924
timestamp 1626908933
transform 1 0 5300 0 1 15318
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1811
timestamp 1626908933
transform 1 0 5136 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3778
timestamp 1626908933
transform 1 0 5136 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1804
timestamp 1626908933
transform 1 0 5136 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3739
timestamp 1626908933
transform 1 0 5136 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1418
timestamp 1626908933
transform 1 0 5520 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3353
timestamp 1626908933
transform 1 0 5520 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1101
timestamp 1626908933
transform 1 0 5088 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_503
timestamp 1626908933
transform 1 0 5088 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_64
timestamp 1626908933
transform -1 0 8160 0 1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_18
timestamp 1626908933
transform -1 0 8160 0 1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_8
timestamp 1626908933
transform 1 0 5088 0 -1 15984
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_6
timestamp 1626908933
transform -1 0 4992 0 1 15984
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_3
timestamp 1626908933
transform 1 0 5088 0 -1 15984
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_1
timestamp 1626908933
transform -1 0 4992 0 1 15984
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_1364
timestamp 1626908933
transform 1 0 6864 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3331
timestamp 1626908933
transform 1 0 6864 0 1 15429
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1447
timestamp 1626908933
transform 1 0 6864 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3382
timestamp 1626908933
transform 1 0 6864 0 1 15429
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1338
timestamp 1626908933
transform 1 0 5616 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3305
timestamp 1626908933
transform 1 0 5616 0 1 15651
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_588
timestamp 1626908933
transform 1 0 6500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1236
timestamp 1626908933
transform 1 0 6500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_588
timestamp 1626908933
transform 1 0 6500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1236
timestamp 1626908933
transform 1 0 6500 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_474
timestamp 1626908933
transform 1 0 7104 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1072
timestamp 1626908933
transform 1 0 7104 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_338
timestamp 1626908933
transform 1 0 7008 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1329
timestamp 1626908933
transform 1 0 7008 0 -1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3603
timestamp 1626908933
transform 1 0 7536 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1636
timestamp 1626908933
transform 1 0 7536 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_544
timestamp 1626908933
transform 1 0 7488 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_187
timestamp 1626908933
transform 1 0 7488 0 -1 15984
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_900
timestamp 1626908933
transform 1 0 7700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_252
timestamp 1626908933
transform 1 0 7700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_900
timestamp 1626908933
transform 1 0 7700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_252
timestamp 1626908933
transform 1 0 7700 0 1 15318
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3577
timestamp 1626908933
transform 1 0 7632 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1642
timestamp 1626908933
transform 1 0 7632 0 1 15725
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3714
timestamp 1626908933
transform 1 0 7824 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1747
timestamp 1626908933
transform 1 0 7824 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_494
timestamp 1626908933
transform 1 0 8160 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1095
timestamp 1626908933
transform 1 0 8160 0 1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1717
timestamp 1626908933
transform 1 0 8016 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3652
timestamp 1626908933
transform 1 0 8016 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_88
timestamp 1626908933
transform 1 0 7584 0 -1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_42
timestamp 1626908933
transform 1 0 7584 0 -1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_39
timestamp 1626908933
transform -1 0 8640 0 1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_100
timestamp 1626908933
transform -1 0 8640 0 1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_33
timestamp 1626908933
transform 1 0 8640 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_85
timestamp 1626908933
transform 1 0 8640 0 1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1736
timestamp 1626908933
transform 1 0 8304 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3703
timestamp 1626908933
transform 1 0 8304 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_495
timestamp 1626908933
transform 1 0 9024 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1096
timestamp 1626908933
transform 1 0 9024 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_48
timestamp 1626908933
transform -1 0 9600 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_110
timestamp 1626908933
transform -1 0 9600 0 1 15984
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_564
timestamp 1626908933
transform 1 0 8900 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1212
timestamp 1626908933
transform 1 0 8900 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_564
timestamp 1626908933
transform 1 0 8900 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1212
timestamp 1626908933
transform 1 0 8900 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_433
timestamp 1626908933
transform 1 0 9600 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1031
timestamp 1626908933
transform 1 0 9600 0 1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1553
timestamp 1626908933
transform 1 0 9264 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3520
timestamp 1626908933
transform 1 0 9264 0 1 15725
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2234
timestamp 1626908933
transform 1 0 9936 0 1 15873
box -29 -23 29 23
use L1M1_PR  L1M1_PR_299
timestamp 1626908933
transform 1 0 9936 0 1 15873
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2245
timestamp 1626908933
transform 1 0 9840 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_278
timestamp 1626908933
transform 1 0 9840 0 1 15873
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_876
timestamp 1626908933
transform 1 0 10100 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_228
timestamp 1626908933
transform 1 0 10100 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_876
timestamp 1626908933
transform 1 0 10100 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_228
timestamp 1626908933
transform 1 0 10100 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_536
timestamp 1626908933
transform 1 0 9984 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_179
timestamp 1626908933
transform 1 0 9984 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_776
timestamp 1626908933
transform 1 0 10272 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_175
timestamp 1626908933
transform 1 0 10272 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_514
timestamp 1626908933
transform 1 0 10464 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1236
timestamp 1626908933
transform 1 0 10464 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_76
timestamp 1626908933
transform -1 0 12768 0 1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_30
timestamp 1626908933
transform -1 0 12768 0 1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_394
timestamp 1626908933
transform 1 0 11328 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_992
timestamp 1626908933
transform 1 0 11328 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_337
timestamp 1626908933
transform 1 0 11232 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1328
timestamp 1626908933
transform 1 0 11232 0 -1 15984
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_540
timestamp 1626908933
transform 1 0 11300 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1188
timestamp 1626908933
transform 1 0 11300 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_540
timestamp 1626908933
transform 1 0 11300 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1188
timestamp 1626908933
transform 1 0 11300 0 1 15984
box -100 -49 100 49
use M1M2_PR  M1M2_PR_59
timestamp 1626908933
transform 1 0 12240 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1460
timestamp 1626908933
transform 1 0 12144 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2026
timestamp 1626908933
transform 1 0 12240 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3427
timestamp 1626908933
transform 1 0 12144 0 1 15577
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_204
timestamp 1626908933
transform 1 0 12500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_852
timestamp 1626908933
transform 1 0 12500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_204
timestamp 1626908933
transform 1 0 12500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_852
timestamp 1626908933
transform 1 0 12500 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_484
timestamp 1626908933
transform 1 0 11712 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1206
timestamp 1626908933
transform 1 0 11712 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_186
timestamp 1626908933
transform 1 0 12480 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_543
timestamp 1626908933
transform 1 0 12480 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_363
timestamp 1626908933
transform 1 0 12768 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_961
timestamp 1626908933
transform 1 0 12768 0 1 15984
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1545
timestamp 1626908933
transform 1 0 12624 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3480
timestamp 1626908933
transform 1 0 12624 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3686
timestamp 1626908933
transform 1 0 13008 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1751
timestamp 1626908933
transform 1 0 13008 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3777
timestamp 1626908933
transform 1 0 13104 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3635
timestamp 1626908933
transform 1 0 13008 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1810
timestamp 1626908933
transform 1 0 13104 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1668
timestamp 1626908933
transform 1 0 13008 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3691
timestamp 1626908933
transform 1 0 13200 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1724
timestamp 1626908933
transform 1 0 13200 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1843
timestamp 1626908933
transform 1 0 13152 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_852
timestamp 1626908933
transform 1 0 13152 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_90
timestamp 1626908933
transform 1 0 13248 0 1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_29
timestamp 1626908933
transform 1 0 13248 0 1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_34
timestamp 1626908933
transform 1 0 13536 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_86
timestamp 1626908933
transform 1 0 13536 0 1 15984
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_516
timestamp 1626908933
transform 1 0 13700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1164
timestamp 1626908933
transform 1 0 13700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_516
timestamp 1626908933
transform 1 0 13700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1164
timestamp 1626908933
transform 1 0 13700 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_68
timestamp 1626908933
transform 1 0 12576 0 -1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_22
timestamp 1626908933
transform 1 0 12576 0 -1 15984
box -38 -49 2726 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_496
timestamp 1626908933
transform 1 0 13920 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1097
timestamp 1626908933
transform 1 0 13920 0 1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_149
timestamp 1626908933
transform 1 0 14064 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2116
timestamp 1626908933
transform 1 0 14064 0 1 15873
box -32 -32 32 32
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_17
timestamp 1626908933
transform -1 0 14688 0 1 15984
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_56
timestamp 1626908933
transform -1 0 14688 0 1 15984
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1098
timestamp 1626908933
transform 1 0 14688 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_497
timestamp 1626908933
transform 1 0 14688 0 1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_67
timestamp 1626908933
transform 1 0 14832 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2002
timestamp 1626908933
transform 1 0 14832 0 1 15429
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_180
timestamp 1626908933
transform 1 0 14900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_828
timestamp 1626908933
transform 1 0 14900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_180
timestamp 1626908933
transform 1 0 14900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_828
timestamp 1626908933
transform 1 0 14900 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_178
timestamp 1626908933
transform 1 0 14976 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_535
timestamp 1626908933
transform 1 0 14976 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_853
timestamp 1626908933
transform 1 0 14880 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1844
timestamp 1626908933
transform 1 0 14880 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3632
timestamp 1626908933
transform 1 0 15120 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1665
timestamp 1626908933
transform 1 0 15120 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1099
timestamp 1626908933
transform 1 0 15072 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_498
timestamp 1626908933
transform 1 0 15072 0 1 15984
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1140
timestamp 1626908933
transform 1 0 16100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_492
timestamp 1626908933
transform 1 0 16100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1140
timestamp 1626908933
transform 1 0 16100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_492
timestamp 1626908933
transform 1 0 16100 0 1 15984
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2099
timestamp 1626908933
transform 1 0 15312 0 1 15873
box -29 -23 29 23
use L1M1_PR  L1M1_PR_164
timestamp 1626908933
transform 1 0 15312 0 1 15873
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2714
timestamp 1626908933
transform 1 0 16560 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_747
timestamp 1626908933
transform 1 0 16560 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_35
timestamp 1626908933
transform -1 0 17568 0 1 15984
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_11
timestamp 1626908933
transform -1 0 17568 0 1 15984
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_36
timestamp 1626908933
transform -1 0 17472 0 -1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_11
timestamp 1626908933
transform -1 0 17472 0 -1 15984
box -38 -49 2246 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_156
timestamp 1626908933
transform 1 0 17300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_804
timestamp 1626908933
transform 1 0 17300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_156
timestamp 1626908933
transform 1 0 17300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_804
timestamp 1626908933
transform 1 0 17300 0 1 15318
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1707
timestamp 1626908933
transform 1 0 16944 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3674
timestamp 1626908933
transform 1 0 16944 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1663
timestamp 1626908933
transform 1 0 17136 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3630
timestamp 1626908933
transform 1 0 17136 0 1 15725
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1746
timestamp 1626908933
transform 1 0 17136 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3681
timestamp 1626908933
transform 1 0 17136 0 1 15725
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1509
timestamp 1626908933
transform 1 0 17424 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3476
timestamp 1626908933
transform 1 0 17424 0 1 15725
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1595
timestamp 1626908933
transform 1 0 17424 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3530
timestamp 1626908933
transform 1 0 17424 0 1 15725
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2815
timestamp 1626908933
transform 1 0 17520 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2814
timestamp 1626908933
transform 1 0 17520 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_848
timestamp 1626908933
transform 1 0 17520 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_847
timestamp 1626908933
transform 1 0 17520 0 1 15725
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1322
timestamp 1626908933
transform 1 0 17568 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_331
timestamp 1626908933
transform 1 0 17568 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_542
timestamp 1626908933
transform 1 0 17472 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_185
timestamp 1626908933
transform 1 0 17472 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2827
timestamp 1626908933
transform 1 0 17616 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2708
timestamp 1626908933
transform 1 0 17712 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_892
timestamp 1626908933
transform 1 0 17616 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_773
timestamp 1626908933
transform 1 0 17712 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3478
timestamp 1626908933
transform 1 0 17808 0 1 15873
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1543
timestamp 1626908933
transform 1 0 17808 0 1 15873
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3426
timestamp 1626908933
transform 1 0 17808 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1459
timestamp 1626908933
transform 1 0 17808 0 1 15873
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2833
timestamp 1626908933
transform 1 0 17904 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2707
timestamp 1626908933
transform 1 0 18000 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_898
timestamp 1626908933
transform 1 0 17904 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_772
timestamp 1626908933
transform 1 0 18000 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1321
timestamp 1626908933
transform 1 0 18048 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_330
timestamp 1626908933
transform 1 0 18048 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2832
timestamp 1626908933
transform 1 0 18096 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2826
timestamp 1626908933
transform 1 0 18192 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_897
timestamp 1626908933
transform 1 0 18096 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_891
timestamp 1626908933
transform 1 0 18192 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1845
timestamp 1626908933
transform 1 0 18144 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_854
timestamp 1626908933
transform 1 0 18144 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_83
timestamp 1626908933
transform 1 0 17952 0 -1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_21
timestamp 1626908933
transform 1 0 17952 0 -1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_77
timestamp 1626908933
transform 1 0 18240 0 -1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_16
timestamp 1626908933
transform 1 0 18240 0 -1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_267
timestamp 1626908933
transform 1 0 17664 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_865
timestamp 1626908933
transform 1 0 17664 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_19
timestamp 1626908933
transform 1 0 17568 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_81
timestamp 1626908933
transform 1 0 17568 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_6
timestamp 1626908933
transform 1 0 18240 0 1 15984
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_45
timestamp 1626908933
transform 1 0 18240 0 1 15984
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2014
timestamp 1626908933
transform 1 0 18576 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_79
timestamp 1626908933
transform 1 0 18576 0 1 15429
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2820
timestamp 1626908933
transform 1 0 18672 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2038
timestamp 1626908933
transform 1 0 18672 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_853
timestamp 1626908933
transform 1 0 18672 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_71
timestamp 1626908933
transform 1 0 18672 0 1 15429
box -32 -32 32 32
use L1M1_PR  L1M1_PR_896
timestamp 1626908933
transform 1 0 18288 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2831
timestamp 1626908933
transform 1 0 18288 0 1 15725
box -29 -23 29 23
use M1M2_PR  M1M2_PR_858
timestamp 1626908933
transform 1 0 18288 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2825
timestamp 1626908933
transform 1 0 18288 0 1 15873
box -32 -32 32 32
use L1M1_PR  L1M1_PR_902
timestamp 1626908933
transform 1 0 18480 0 1 15873
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2837
timestamp 1626908933
transform 1 0 18480 0 1 15873
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_468
timestamp 1626908933
transform 1 0 18500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1116
timestamp 1626908933
transform 1 0 18500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_468
timestamp 1626908933
transform 1 0 18500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1116
timestamp 1626908933
transform 1 0 18500 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_775
timestamp 1626908933
transform 1 0 18528 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_174
timestamp 1626908933
transform 1 0 18528 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_12
timestamp 1626908933
transform 1 0 19104 0 -1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_74
timestamp 1626908933
transform 1 0 19104 0 -1 15984
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_244
timestamp 1626908933
transform 1 0 18720 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_842
timestamp 1626908933
transform 1 0 18720 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_5
timestamp 1626908933
transform 1 0 18816 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_57
timestamp 1626908933
transform 1 0 18816 0 1 15984
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2627
timestamp 1626908933
transform 1 0 19248 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_692
timestamp 1626908933
transform 1 0 19248 0 1 15429
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2640
timestamp 1626908933
transform 1 0 19248 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_673
timestamp 1626908933
transform 1 0 19248 0 1 15429
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2019
timestamp 1626908933
transform 1 0 19152 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_84
timestamp 1626908933
transform 1 0 19152 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2717
timestamp 1626908933
transform 1 0 19344 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_782
timestamp 1626908933
transform 1 0 19344 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2721
timestamp 1626908933
transform 1 0 19344 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_754
timestamp 1626908933
transform 1 0 19344 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_326
timestamp 1626908933
transform 1 0 19200 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1048
timestamp 1626908933
transform 1 0 19200 0 1 15984
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_780
timestamp 1626908933
transform 1 0 19700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_132
timestamp 1626908933
transform 1 0 19700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_780
timestamp 1626908933
transform 1 0 19700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_132
timestamp 1626908933
transform 1 0 19700 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1327
timestamp 1626908933
transform 1 0 19392 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_336
timestamp 1626908933
transform 1 0 19392 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2017
timestamp 1626908933
transform 1 0 20016 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_82
timestamp 1626908933
transform 1 0 20016 0 1 15577
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2040
timestamp 1626908933
transform 1 0 19920 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_73
timestamp 1626908933
transform 1 0 19920 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1326
timestamp 1626908933
transform 1 0 19872 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_335
timestamp 1626908933
transform 1 0 19872 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_534
timestamp 1626908933
transform 1 0 19968 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_177
timestamp 1626908933
transform 1 0 19968 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_827
timestamp 1626908933
transform 1 0 19488 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_229
timestamp 1626908933
transform 1 0 19488 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_329
timestamp 1626908933
transform 1 0 20448 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1320
timestamp 1626908933
transform 1 0 20448 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_854
timestamp 1626908933
transform 1 0 20112 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1693
timestamp 1626908933
transform 1 0 20592 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2821
timestamp 1626908933
transform 1 0 20112 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3660
timestamp 1626908933
transform 1 0 20592 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_32
timestamp 1626908933
transform 1 0 20064 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_94
timestamp 1626908933
transform 1 0 20064 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_300
timestamp 1626908933
transform 1 0 20544 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1022
timestamp 1626908933
transform 1 0 20544 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_19
timestamp 1626908933
transform -1 0 21888 0 1 15984
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_58
timestamp 1626908933
transform -1 0 21888 0 1 15984
box -38 -49 614 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_444
timestamp 1626908933
transform 1 0 20900 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1092
timestamp 1626908933
transform 1 0 20900 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_444
timestamp 1626908933
transform 1 0 20900 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1092
timestamp 1626908933
transform 1 0 20900 0 1 15984
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3623
timestamp 1626908933
transform 1 0 21552 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1656
timestamp 1626908933
transform 1 0 21552 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3676
timestamp 1626908933
transform 1 0 21840 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1741
timestamp 1626908933
transform 1 0 21840 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3421
timestamp 1626908933
transform 1 0 21936 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1454
timestamp 1626908933
transform 1 0 21936 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1319
timestamp 1626908933
transform 1 0 21888 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_328
timestamp 1626908933
transform 1 0 21888 0 1 15984
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_756
timestamp 1626908933
transform 1 0 22100 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_108
timestamp 1626908933
transform 1 0 22100 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_756
timestamp 1626908933
transform 1 0 22100 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_108
timestamp 1626908933
transform 1 0 22100 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_273
timestamp 1626908933
transform 1 0 21984 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_995
timestamp 1626908933
transform 1 0 21984 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_37
timestamp 1626908933
transform -1 0 22272 0 -1 15984
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_13
timestamp 1626908933
transform -1 0 22272 0 -1 15984
box -38 -49 2342 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_184
timestamp 1626908933
transform 1 0 22464 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_541
timestamp 1626908933
transform 1 0 22464 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_490
timestamp 1626908933
transform 1 0 22272 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1091
timestamp 1626908933
transform 1 0 22272 0 -1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1539
timestamp 1626908933
transform 1 0 22224 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3474
timestamp 1626908933
transform 1 0 22224 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_327
timestamp 1626908933
transform 1 0 22752 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1318
timestamp 1626908933
transform 1 0 22752 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_249
timestamp 1626908933
transform 1 0 22560 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_971
timestamp 1626908933
transform 1 0 22560 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_173
timestamp 1626908933
transform 1 0 22848 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_771
timestamp 1626908933
transform 1 0 22848 0 1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3657
timestamp 1626908933
transform 1 0 22992 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1690
timestamp 1626908933
transform 1 0 22992 0 1 15503
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1068
timestamp 1626908933
transform 1 0 23300 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_420
timestamp 1626908933
transform 1 0 23300 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1068
timestamp 1626908933
transform 1 0 23300 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_420
timestamp 1626908933
transform 1 0 23300 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_774
timestamp 1626908933
transform 1 0 23328 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_770
timestamp 1626908933
transform 1 0 23232 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_173
timestamp 1626908933
transform 1 0 23328 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_169
timestamp 1626908933
transform 1 0 23232 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_159
timestamp 1626908933
transform 1 0 23520 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_757
timestamp 1626908933
transform 1 0 23520 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_2
timestamp 1626908933
transform 1 0 23424 0 1 15984
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_17
timestamp 1626908933
transform 1 0 23424 0 1 15984
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_326
timestamp 1626908933
transform 1 0 24096 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1317
timestamp 1626908933
transform 1 0 24096 0 1 15984
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_84
timestamp 1626908933
transform 1 0 24500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_732
timestamp 1626908933
transform 1 0 24500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_84
timestamp 1626908933
transform 1 0 24500 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_732
timestamp 1626908933
transform 1 0 24500 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_203
timestamp 1626908933
transform 1 0 24192 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_219
timestamp 1626908933
transform 1 0 23904 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_925
timestamp 1626908933
transform 1 0 24192 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_941
timestamp 1626908933
transform 1 0 23904 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1325
timestamp 1626908933
transform 1 0 24672 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_334
timestamp 1626908933
transform 1 0 24672 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_731
timestamp 1626908933
transform 1 0 24768 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_133
timestamp 1626908933
transform 1 0 24768 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_176
timestamp 1626908933
transform 1 0 24960 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_533
timestamp 1626908933
transform 1 0 24960 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_325
timestamp 1626908933
transform 1 0 25056 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1316
timestamp 1626908933
transform 1 0 25056 0 1 15984
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_396
timestamp 1626908933
transform 1 0 25700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1044
timestamp 1626908933
transform 1 0 25700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_396
timestamp 1626908933
transform 1 0 25700 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1044
timestamp 1626908933
transform 1 0 25700 0 1 15984
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_185
timestamp 1626908933
transform 1 0 25152 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_186
timestamp 1626908933
transform 1 0 25152 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_907
timestamp 1626908933
transform 1 0 25152 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_908
timestamp 1626908933
transform 1 0 25152 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_172
timestamp 1626908933
transform 1 0 25920 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_773
timestamp 1626908933
transform 1 0 25920 0 -1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1419
timestamp 1626908933
transform 1 0 26256 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1895
timestamp 1626908933
transform 1 0 26352 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3386
timestamp 1626908933
transform 1 0 26256 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3862
timestamp 1626908933
transform 1 0 26352 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_156
timestamp 1626908933
transform 1 0 26496 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_878
timestamp 1626908933
transform 1 0 26496 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_105
timestamp 1626908933
transform 1 0 26112 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_703
timestamp 1626908933
transform 1 0 26112 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_3
timestamp 1626908933
transform 1 0 25920 0 1 15984
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_18
timestamp 1626908933
transform 1 0 25920 0 1 15984
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_324
timestamp 1626908933
transform 1 0 26976 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1315
timestamp 1626908933
transform 1 0 26976 0 1 15984
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_60
timestamp 1626908933
transform 1 0 26900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_708
timestamp 1626908933
transform 1 0 26900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_60
timestamp 1626908933
transform 1 0 26900 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_708
timestamp 1626908933
transform 1 0 26900 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_333
timestamp 1626908933
transform 1 0 27264 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_849
timestamp 1626908933
transform 1 0 27360 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1324
timestamp 1626908933
transform 1 0 27264 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1840
timestamp 1626908933
transform 1 0 27360 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_141
timestamp 1626908933
transform 1 0 27072 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_863
timestamp 1626908933
transform 1 0 27072 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_94
timestamp 1626908933
transform 1 0 26592 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_692
timestamp 1626908933
transform 1 0 26592 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_772
timestamp 1626908933
transform 1 0 27552 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_171
timestamp 1626908933
transform 1 0 27552 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_540
timestamp 1626908933
transform 1 0 27456 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_183
timestamp 1626908933
transform 1 0 27456 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_168
timestamp 1626908933
transform 1 0 27840 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_769
timestamp 1626908933
transform 1 0 27840 0 1 15984
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_372
timestamp 1626908933
transform 1 0 28100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1020
timestamp 1626908933
transform 1 0 28100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_372
timestamp 1626908933
transform 1 0 28100 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1020
timestamp 1626908933
transform 1 0 28100 0 1 15984
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1347
timestamp 1626908933
transform 1 0 28272 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1402
timestamp 1626908933
transform 1 0 28464 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3314
timestamp 1626908933
transform 1 0 28272 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3369
timestamp 1626908933
transform 1 0 28464 0 1 15429
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1428
timestamp 1626908933
transform 1 0 28176 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1505
timestamp 1626908933
transform 1 0 28368 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3363
timestamp 1626908933
transform 1 0 28176 0 1 15725
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3440
timestamp 1626908933
transform 1 0 28368 0 1 15725
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_107
timestamp 1626908933
transform 1 0 28416 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_829
timestamp 1626908933
transform 1 0 28416 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_74
timestamp 1626908933
transform 1 0 28032 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_78
timestamp 1626908933
transform 1 0 27744 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_672
timestamp 1626908933
transform 1 0 28032 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_676
timestamp 1626908933
transform 1 0 27744 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_12
timestamp 1626908933
transform 1 0 28128 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_37
timestamp 1626908933
transform 1 0 28128 0 -1 15984
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1485
timestamp 1626908933
transform 1 0 28560 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3420
timestamp 1626908933
transform 1 0 28560 0 1 15429
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_36
timestamp 1626908933
transform 1 0 29300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_684
timestamp 1626908933
transform 1 0 29300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_36
timestamp 1626908933
transform 1 0 29300 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_684
timestamp 1626908933
transform 1 0 29300 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_74
timestamp 1626908933
transform 1 0 29184 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_91
timestamp 1626908933
transform 1 0 28992 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_796
timestamp 1626908933
transform 1 0 29184 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_813
timestamp 1626908933
transform 1 0 28992 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_49
timestamp 1626908933
transform 1 0 28608 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_647
timestamp 1626908933
transform 1 0 28608 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_491
timestamp 1626908933
transform 1 0 29760 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1092
timestamp 1626908933
transform 1 0 29760 0 -1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_414
timestamp 1626908933
transform 1 0 29424 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2381
timestamp 1626908933
transform 1 0 29424 0 1 15725
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2326
timestamp 1626908933
transform 1 0 29904 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_359
timestamp 1626908933
transform 1 0 29904 0 1 15873
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_532
timestamp 1626908933
transform 1 0 29952 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_175
timestamp 1626908933
transform 1 0 29952 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3752
timestamp 1626908933
transform 1 0 30096 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2317
timestamp 1626908933
transform 1 0 30000 0 1 15873
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1817
timestamp 1626908933
transform 1 0 30096 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_382
timestamp 1626908933
transform 1 0 30000 0 1 15873
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3797
timestamp 1626908933
transform 1 0 30096 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1830
timestamp 1626908933
transform 1 0 30096 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_768
timestamp 1626908933
transform 1 0 30048 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_167
timestamp 1626908933
transform 1 0 30048 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_4
timestamp 1626908933
transform 1 0 29952 0 -1 15984
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_19
timestamp 1626908933
transform 1 0 29952 0 -1 15984
box -38 -49 710 715
use L1M1_PR  L1M1_PR_3796
timestamp 1626908933
transform 1 0 30384 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2343
timestamp 1626908933
transform 1 0 30288 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1861
timestamp 1626908933
transform 1 0 30384 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_408
timestamp 1626908933
transform 1 0 30288 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1314
timestamp 1626908933
transform 1 0 30240 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_323
timestamp 1626908933
transform 1 0 30240 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_768
timestamp 1626908933
transform 1 0 30336 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_46
timestamp 1626908933
transform 1 0 30336 0 1 15984
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_996
timestamp 1626908933
transform 1 0 30500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_348
timestamp 1626908933
transform 1 0 30500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_996
timestamp 1626908933
transform 1 0 30500 0 1 15984
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_348
timestamp 1626908933
transform 1 0 30500 0 1 15984
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3733
timestamp 1626908933
transform 1 0 30576 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1798
timestamp 1626908933
transform 1 0 30576 0 1 15429
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3852
timestamp 1626908933
transform 1 0 30672 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1885
timestamp 1626908933
transform 1 0 30672 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1323
timestamp 1626908933
transform 1 0 30816 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_332
timestamp 1626908933
transform 1 0 30816 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_771
timestamp 1626908933
transform 1 0 30624 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_170
timestamp 1626908933
transform 1 0 30624 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_322
timestamp 1626908933
transform 1 0 31104 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1313
timestamp 1626908933
transform 1 0 31104 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1794
timestamp 1626908933
transform 1 0 30960 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3761
timestamp 1626908933
transform 1 0 30960 0 1 15429
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_11
timestamp 1626908933
transform 1 0 31200 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_28
timestamp 1626908933
transform 1 0 30912 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_733
timestamp 1626908933
transform 1 0 31200 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_750
timestamp 1626908933
transform 1 0 30912 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_182
timestamp 1626908933
transform 1 0 31680 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_539
timestamp 1626908933
transform 1 0 31680 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_492
timestamp 1626908933
transform 1 0 31776 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1093
timestamp 1626908933
transform 1 0 31776 0 -1 15984
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_12
timestamp 1626908933
transform 1 0 31700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_660
timestamp 1626908933
transform 1 0 31700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_12
timestamp 1626908933
transform 1 0 31700 0 1 15318
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_660
timestamp 1626908933
transform 1 0 31700 0 1 15318
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_850
timestamp 1626908933
transform 1 0 31968 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_855
timestamp 1626908933
transform 1 0 31968 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1841
timestamp 1626908933
transform 1 0 31968 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1846
timestamp 1626908933
transform 1 0 31968 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_166
timestamp 1626908933
transform 1 0 0 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_767
timestamp 1626908933
transform 1 0 0 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1880
timestamp 1626908933
transform 1 0 240 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1947
timestamp 1626908933
transform 1 0 48 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1966
timestamp 1626908933
transform 1 0 48 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3847
timestamp 1626908933
transform 1 0 240 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3914
timestamp 1626908933
transform 1 0 48 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3933
timestamp 1626908933
transform 1 0 48 0 1 16391
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1731
timestamp 1626908933
transform 1 0 816 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3666
timestamp 1626908933
transform 1 0 816 0 1 16539
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_323
timestamp 1626908933
transform 1 0 500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_971
timestamp 1626908933
transform 1 0 500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_323
timestamp 1626908933
transform 1 0 500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_971
timestamp 1626908933
transform 1 0 500 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_711
timestamp 1626908933
transform 1 0 192 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1433
timestamp 1626908933
transform 1 0 192 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1312
timestamp 1626908933
transform 1 0 960 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_321
timestamp 1626908933
transform 1 0 960 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1171
timestamp 1626908933
transform 1 0 1056 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_573
timestamp 1626908933
transform 1 0 1056 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1399
timestamp 1626908933
transform 1 0 1440 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_677
timestamp 1626908933
transform 1 0 1440 0 -1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3930
timestamp 1626908933
transform 1 0 2448 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1963
timestamp 1626908933
transform 1 0 2448 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1311
timestamp 1626908933
transform 1 0 2208 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_320
timestamp 1626908933
transform 1 0 2208 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1100
timestamp 1626908933
transform 1 0 2304 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_499
timestamp 1626908933
transform 1 0 2304 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_531
timestamp 1626908933
transform 1 0 2496 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_174
timestamp 1626908933
transform 1 0 2496 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3868
timestamp 1626908933
transform 1 0 2640 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1933
timestamp 1626908933
transform 1 0 2640 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3615
timestamp 1626908933
transform 1 0 2736 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1648
timestamp 1626908933
transform 1 0 2736 0 1 16539
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_87
timestamp 1626908933
transform 1 0 2592 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_35
timestamp 1626908933
transform 1 0 2592 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_856
timestamp 1626908933
transform 1 0 2976 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1847
timestamp 1626908933
transform 1 0 2976 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1916
timestamp 1626908933
transform 1 0 3024 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3851
timestamp 1626908933
transform 1 0 3024 0 1 16243
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_299
timestamp 1626908933
transform 1 0 2900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_947
timestamp 1626908933
transform 1 0 2900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_299
timestamp 1626908933
transform 1 0 2900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_947
timestamp 1626908933
transform 1 0 2900 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_319
timestamp 1626908933
transform 1 0 3456 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1310
timestamp 1626908933
transform 1 0 3456 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1602
timestamp 1626908933
transform 1 0 3408 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3569
timestamp 1626908933
transform 1 0 3408 0 1 16095
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1695
timestamp 1626908933
transform 1 0 3408 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3630
timestamp 1626908933
transform 1 0 3408 0 1 16095
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_628
timestamp 1626908933
transform 1 0 3552 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1350
timestamp 1626908933
transform 1 0 3552 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_49
timestamp 1626908933
transform -1 0 3456 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_111
timestamp 1626908933
transform -1 0 3456 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_104
timestamp 1626908933
transform 1 0 4320 0 -1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_42
timestamp 1626908933
transform 1 0 4320 0 -1 17316
box -38 -49 326 715
use M1M2_PR  M1M2_PR_402
timestamp 1626908933
transform 1 0 4656 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2369
timestamp 1626908933
transform 1 0 4656 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_400
timestamp 1626908933
transform 1 0 4560 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1915
timestamp 1626908933
transform 1 0 4944 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2335
timestamp 1626908933
transform 1 0 4560 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3850
timestamp 1626908933
transform 1 0 4944 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1106
timestamp 1626908933
transform 1 0 4848 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3073
timestamp 1626908933
transform 1 0 4848 0 1 16539
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_275
timestamp 1626908933
transform 1 0 5300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_923
timestamp 1626908933
transform 1 0 5300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_275
timestamp 1626908933
transform 1 0 5300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_923
timestamp 1626908933
transform 1 0 5300 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_621
timestamp 1626908933
transform 1 0 4608 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1343
timestamp 1626908933
transform 1 0 4608 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_1
timestamp 1626908933
transform 1 0 5376 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_70
timestamp 1626908933
transform 1 0 5376 0 -1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2239
timestamp 1626908933
transform 1 0 5808 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_304
timestamp 1626908933
transform 1 0 5808 0 1 16169
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1089
timestamp 1626908933
transform 1 0 5856 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_491
timestamp 1626908933
transform 1 0 5856 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1101
timestamp 1626908933
transform 1 0 6720 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_500
timestamp 1626908933
transform 1 0 6720 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_3
timestamp 1626908933
transform 1 0 6240 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_0
timestamp 1626908933
transform 1 0 6240 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_44
timestamp 1626908933
transform 1 0 7008 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_19
timestamp 1626908933
transform 1 0 7008 0 -1 17316
box -38 -49 518 715
use M1M2_PR  M1M2_PR_3912
timestamp 1626908933
transform 1 0 7248 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1945
timestamp 1626908933
transform 1 0 7248 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1848
timestamp 1626908933
transform 1 0 6912 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_857
timestamp 1626908933
transform 1 0 6912 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_530
timestamp 1626908933
transform 1 0 7488 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_173
timestamp 1626908933
transform 1 0 7488 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1635
timestamp 1626908933
transform 1 0 7536 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3602
timestamp 1626908933
transform 1 0 7536 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1720
timestamp 1626908933
transform 1 0 7728 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3655
timestamp 1626908933
transform 1 0 7728 0 1 16317
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_251
timestamp 1626908933
transform 1 0 7700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_899
timestamp 1626908933
transform 1 0 7700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_251
timestamp 1626908933
transform 1 0 7700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_899
timestamp 1626908933
transform 1 0 7700 0 1 16650
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3575
timestamp 1626908933
transform 1 0 8112 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1640
timestamp 1626908933
transform 1 0 8112 0 1 16391
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3713
timestamp 1626908933
transform 1 0 7824 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3518
timestamp 1626908933
transform 1 0 8112 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1746
timestamp 1626908933
transform 1 0 7824 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1551
timestamp 1626908933
transform 1 0 8112 0 1 16391
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3574
timestamp 1626908933
transform 1 0 8112 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1639
timestamp 1626908933
transform 1 0 8112 0 1 16761
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3517
timestamp 1626908933
transform 1 0 8112 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1550
timestamp 1626908933
transform 1 0 8112 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1849
timestamp 1626908933
transform 1 0 7968 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_858
timestamp 1626908933
transform 1 0 7968 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_467
timestamp 1626908933
transform 1 0 7584 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1065
timestamp 1626908933
transform 1 0 7584 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_35
timestamp 1626908933
transform 1 0 8064 0 -1 17316
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_74
timestamp 1626908933
transform 1 0 8064 0 -1 17316
box -38 -49 614 715
use M1M2_PR  M1M2_PR_281
timestamp 1626908933
transform 1 0 8496 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1104
timestamp 1626908933
transform 1 0 8400 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2248
timestamp 1626908933
transform 1 0 8496 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3071
timestamp 1626908933
transform 1 0 8400 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_302
timestamp 1626908933
transform 1 0 8304 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1171
timestamp 1626908933
transform 1 0 8496 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2237
timestamp 1626908933
transform 1 0 8304 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3106
timestamp 1626908933
transform 1 0 8496 0 1 16539
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_501
timestamp 1626908933
transform 1 0 8640 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1102
timestamp 1626908933
transform 1 0 8640 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_859
timestamp 1626908933
transform 1 0 8832 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1850
timestamp 1626908933
transform 1 0 8832 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1732
timestamp 1626908933
transform 1 0 8688 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3699
timestamp 1626908933
transform 1 0 8688 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1102
timestamp 1626908933
transform 1 0 9072 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3069
timestamp 1626908933
transform 1 0 9072 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1169
timestamp 1626908933
transform 1 0 9072 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3104
timestamp 1626908933
transform 1 0 9072 0 1 16539
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_502
timestamp 1626908933
transform 1 0 9216 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1103
timestamp 1626908933
transform 1 0 9216 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1098
timestamp 1626908933
transform 1 0 9264 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1552
timestamp 1626908933
transform 1 0 9264 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3065
timestamp 1626908933
transform 1 0 9264 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3519
timestamp 1626908933
transform 1 0 9264 0 1 16095
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1641
timestamp 1626908933
transform 1 0 9360 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3576
timestamp 1626908933
transform 1 0 9360 0 1 16095
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_120
timestamp 1626908933
transform -1 0 9888 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_51
timestamp 1626908933
transform -1 0 9888 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_43
timestamp 1626908933
transform 1 0 8928 0 -1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_105
timestamp 1626908933
transform 1 0 8928 0 -1 17316
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1100
timestamp 1626908933
transform 1 0 9456 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3067
timestamp 1626908933
transform 1 0 9456 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1162
timestamp 1626908933
transform 1 0 9552 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1166
timestamp 1626908933
transform 1 0 9456 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3097
timestamp 1626908933
transform 1 0 9552 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3101
timestamp 1626908933
transform 1 0 9456 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_503
timestamp 1626908933
transform 1 0 9888 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1104
timestamp 1626908933
transform 1 0 9888 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_277
timestamp 1626908933
transform 1 0 9840 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2244
timestamp 1626908933
transform 1 0 9840 0 1 16761
box -32 -32 32 32
use L1M1_PR  L1M1_PR_298
timestamp 1626908933
transform 1 0 9936 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2233
timestamp 1626908933
transform 1 0 9936 0 1 16761
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_860
timestamp 1626908933
transform 1 0 10080 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1851
timestamp 1626908933
transform 1 0 10080 0 -1 17316
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_227
timestamp 1626908933
transform 1 0 10100 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_875
timestamp 1626908933
transform 1 0 10100 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_227
timestamp 1626908933
transform 1 0 10100 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_875
timestamp 1626908933
transform 1 0 10100 0 1 16650
box -100 -49 100 49
use M1M2_PR  M1M2_PR_218
timestamp 1626908933
transform 1 0 10320 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2185
timestamp 1626908933
transform 1 0 10320 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_238
timestamp 1626908933
transform 1 0 10512 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2173
timestamp 1626908933
transform 1 0 10512 0 1 16539
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_112
timestamp 1626908933
transform -1 0 10656 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_43
timestamp 1626908933
transform -1 0 10656 0 -1 17316
box -38 -49 518 715
use M1M2_PR  M1M2_PR_2902
timestamp 1626908933
transform 1 0 10992 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2243
timestamp 1626908933
transform 1 0 10800 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_935
timestamp 1626908933
transform 1 0 10992 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_276
timestamp 1626908933
transform 1 0 10800 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_766
timestamp 1626908933
transform 1 0 10656 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_165
timestamp 1626908933
transform 1 0 10656 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1003
timestamp 1626908933
transform 1 0 10848 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_405
timestamp 1626908933
transform 1 0 10848 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_318
timestamp 1626908933
transform 1 0 11616 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1309
timestamp 1626908933
transform 1 0 11616 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1674
timestamp 1626908933
transform 1 0 11280 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3609
timestamp 1626908933
transform 1 0 11280 0 1 16761
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_40
timestamp 1626908933
transform -1 0 11616 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_102
timestamp 1626908933
transform -1 0 11616 0 -1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1623
timestamp 1626908933
transform 1 0 12336 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3590
timestamp 1626908933
transform 1 0 12336 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1709
timestamp 1626908933
transform 1 0 12336 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3644
timestamp 1626908933
transform 1 0 12336 0 1 16317
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_203
timestamp 1626908933
transform 1 0 12500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_851
timestamp 1626908933
transform 1 0 12500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_203
timestamp 1626908933
transform 1 0 12500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_851
timestamp 1626908933
transform 1 0 12500 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_483
timestamp 1626908933
transform 1 0 11712 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1205
timestamp 1626908933
transform 1 0 11712 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_172
timestamp 1626908933
transform 1 0 12480 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_529
timestamp 1626908933
transform 1 0 12480 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1584
timestamp 1626908933
transform 1 0 12720 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1585
timestamp 1626908933
transform 1 0 12720 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3551
timestamp 1626908933
transform 1 0 12720 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3552
timestamp 1626908933
transform 1 0 12720 0 1 16391
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1673
timestamp 1626908933
transform 1 0 12720 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3608
timestamp 1626908933
transform 1 0 12720 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_991
timestamp 1626908933
transform 1 0 13296 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2926
timestamp 1626908933
transform 1 0 13296 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_167
timestamp 1626908933
transform 1 0 13488 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_997
timestamp 1626908933
transform 1 0 13584 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2102
timestamp 1626908933
transform 1 0 13488 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2932
timestamp 1626908933
transform 1 0 13584 0 1 16243
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_87
timestamp 1626908933
transform -1 0 15264 0 -1 17316
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_41
timestamp 1626908933
transform -1 0 15264 0 -1 17316
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_148
timestamp 1626908933
transform 1 0 14064 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2115
timestamp 1626908933
transform 1 0 14064 0 1 16169
box -32 -32 32 32
use L1M1_PR  L1M1_PR_166
timestamp 1626908933
transform 1 0 14064 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2101
timestamp 1626908933
transform 1 0 14064 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_990
timestamp 1626908933
transform 1 0 14256 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2925
timestamp 1626908933
transform 1 0 14256 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_996
timestamp 1626908933
transform 1 0 14448 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2931
timestamp 1626908933
transform 1 0 14448 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1596
timestamp 1626908933
transform 1 0 14640 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3531
timestamp 1626908933
transform 1 0 14640 0 1 16169
box -29 -23 29 23
use L1M1_PR  L1M1_PR_75
timestamp 1626908933
transform 1 0 15312 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2010
timestamp 1626908933
transform 1 0 15312 0 1 16095
box -29 -23 29 23
use M1M2_PR  M1M2_PR_938
timestamp 1626908933
transform 1 0 15504 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2905
timestamp 1626908933
transform 1 0 15504 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_66
timestamp 1626908933
transform 1 0 16272 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2033
timestamp 1626908933
transform 1 0 16272 0 1 16095
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_827
timestamp 1626908933
transform 1 0 14900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_179
timestamp 1626908933
transform 1 0 14900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_827
timestamp 1626908933
transform 1 0 14900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_179
timestamp 1626908933
transform 1 0 14900 0 1 16650
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2121
timestamp 1626908933
transform 1 0 15888 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_154
timestamp 1626908933
transform 1 0 15888 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_37
timestamp 1626908933
transform 1 0 15264 0 -1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_12
timestamp 1626908933
transform 1 0 15264 0 -1 17316
box -38 -49 2246 715
use M1M2_PR  M1M2_PR_1706
timestamp 1626908933
transform 1 0 16944 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3673
timestamp 1626908933
transform 1 0 16944 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1662
timestamp 1626908933
transform 1 0 17136 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3629
timestamp 1626908933
transform 1 0 17136 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1745
timestamp 1626908933
transform 1 0 17136 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3680
timestamp 1626908933
transform 1 0 17136 0 1 16317
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_155
timestamp 1626908933
transform 1 0 17300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_803
timestamp 1626908933
transform 1 0 17300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_155
timestamp 1626908933
transform 1 0 17300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_803
timestamp 1626908933
transform 1 0 17300 0 1 16650
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3479
timestamp 1626908933
transform 1 0 17520 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1544
timestamp 1626908933
transform 1 0 17520 0 1 16243
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3475
timestamp 1626908933
transform 1 0 17424 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1508
timestamp 1626908933
transform 1 0 17424 0 1 16169
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2105
timestamp 1626908933
transform 1 0 17424 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_170
timestamp 1626908933
transform 1 0 17424 0 1 16761
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1105
timestamp 1626908933
transform 1 0 17568 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_504
timestamp 1626908933
transform 1 0 17568 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_528
timestamp 1626908933
transform 1 0 17472 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_171
timestamp 1626908933
transform 1 0 17472 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_861
timestamp 1626908933
transform 1 0 17760 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1852
timestamp 1626908933
transform 1 0 17760 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1458
timestamp 1626908933
transform 1 0 17808 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3425
timestamp 1626908933
transform 1 0 17808 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_69
timestamp 1626908933
transform 1 0 18768 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2036
timestamp 1626908933
transform 1 0 18768 0 1 16095
box -32 -32 32 32
use L1M1_PR  L1M1_PR_78
timestamp 1626908933
transform 1 0 18864 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2013
timestamp 1626908933
transform 1 0 18864 0 1 16095
box -29 -23 29 23
use M1M2_PR  M1M2_PR_857
timestamp 1626908933
transform 1 0 18288 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2824
timestamp 1626908933
transform 1 0 18288 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_901
timestamp 1626908933
transform 1 0 18480 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2836
timestamp 1626908933
transform 1 0 18480 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_852
timestamp 1626908933
transform 1 0 18672 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2819
timestamp 1626908933
transform 1 0 18672 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_895
timestamp 1626908933
transform 1 0 18672 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2830
timestamp 1626908933
transform 1 0 18672 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_753
timestamp 1626908933
transform 1 0 19344 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2720
timestamp 1626908933
transform 1 0 19344 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1457
timestamp 1626908933
transform 1 0 18192 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3424
timestamp 1626908933
transform 1 0 18192 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1541
timestamp 1626908933
transform 1 0 18288 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3476
timestamp 1626908933
transform 1 0 18288 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_70
timestamp 1626908933
transform 1 0 18672 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2037
timestamp 1626908933
transform 1 0 18672 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_36
timestamp 1626908933
transform 1 0 17856 0 -1 17316
box -38 -49 2342 715
use sky130_fd_sc_hs__dfrbp_1  sky130_fd_sc_hs__dfrbp_1_12
timestamp 1626908933
transform 1 0 17856 0 -1 17316
box -38 -49 2342 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_131
timestamp 1626908933
transform 1 0 19700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_779
timestamp 1626908933
transform 1 0 19700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_131
timestamp 1626908933
transform 1 0 19700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_779
timestamp 1626908933
transform 1 0 19700 0 1 16650
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2936
timestamp 1626908933
transform 1 0 20112 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1001
timestamp 1626908933
transform 1 0 20112 0 1 16243
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2908
timestamp 1626908933
transform 1 0 19920 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_941
timestamp 1626908933
transform 1 0 19920 0 1 16243
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2011
timestamp 1626908933
transform 1 0 20112 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_76
timestamp 1626908933
transform 1 0 20112 0 1 16761
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3470
timestamp 1626908933
transform 1 0 20112 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1503
timestamp 1626908933
transform 1 0 20112 0 1 16539
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_765
timestamp 1626908933
transform 1 0 20160 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_164
timestamp 1626908933
transform 1 0 20160 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_317
timestamp 1626908933
transform 1 0 20352 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1308
timestamp 1626908933
transform 1 0 20352 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_779
timestamp 1626908933
transform 1 0 20208 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1007
timestamp 1626908933
transform 1 0 20400 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1589
timestamp 1626908933
transform 1 0 20400 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2714
timestamp 1626908933
transform 1 0 20208 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2942
timestamp 1626908933
transform 1 0 20400 0 1 16243
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3524
timestamp 1626908933
transform 1 0 20400 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_947
timestamp 1626908933
transform 1 0 20976 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2914
timestamp 1626908933
transform 1 0 20976 0 1 16243
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_299
timestamp 1626908933
transform 1 0 20448 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1021
timestamp 1626908933
transform 1 0 20448 0 -1 17316
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2940
timestamp 1626908933
transform 1 0 21456 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2116
timestamp 1626908933
transform 1 0 21360 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1005
timestamp 1626908933
transform 1 0 21456 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_181
timestamp 1626908933
transform 1 0 21360 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2131
timestamp 1626908933
transform 1 0 21360 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_164
timestamp 1626908933
transform 1 0 21360 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2947
timestamp 1626908933
transform 1 0 21360 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1012
timestamp 1626908933
transform 1 0 21360 0 1 16761
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_88
timestamp 1626908933
transform 1 0 21216 0 -1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_27
timestamp 1626908933
transform 1 0 21216 0 -1 17316
box -38 -49 326 715
use L1M1_PR  L1M1_PR_2946
timestamp 1626908933
transform 1 0 21648 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1011
timestamp 1626908933
transform 1 0 21648 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2918
timestamp 1626908933
transform 1 0 21648 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_951
timestamp 1626908933
transform 1 0 21648 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3523
timestamp 1626908933
transform 1 0 21840 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1588
timestamp 1626908933
transform 1 0 21840 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2917
timestamp 1626908933
transform 1 0 21648 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_950
timestamp 1626908933
transform 1 0 21648 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_764
timestamp 1626908933
transform 1 0 21504 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_163
timestamp 1626908933
transform 1 0 21504 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_272
timestamp 1626908933
transform 1 0 21696 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_994
timestamp 1626908933
transform 1 0 21696 0 -1 17316
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_755
timestamp 1626908933
transform 1 0 22100 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_107
timestamp 1626908933
transform 1 0 22100 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_755
timestamp 1626908933
transform 1 0 22100 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_107
timestamp 1626908933
transform 1 0 22100 0 1 16650
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3801
timestamp 1626908933
transform 1 0 21936 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1834
timestamp 1626908933
transform 1 0 21936 0 1 16391
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3754
timestamp 1626908933
transform 1 0 23376 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2323
timestamp 1626908933
transform 1 0 23472 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1819
timestamp 1626908933
transform 1 0 23376 0 1 16391
box -29 -23 29 23
use L1M1_PR  L1M1_PR_388
timestamp 1626908933
transform 1 0 23472 0 1 16095
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2332
timestamp 1626908933
transform 1 0 22992 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_365
timestamp 1626908933
transform 1 0 22992 0 1 16095
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_527
timestamp 1626908933
transform 1 0 22464 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_170
timestamp 1626908933
transform 1 0 22464 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1501
timestamp 1626908933
transform 1 0 23760 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1899
timestamp 1626908933
transform 1 0 23856 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3468
timestamp 1626908933
transform 1 0 23760 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3866
timestamp 1626908933
transform 1 0 23856 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_414
timestamp 1626908933
transform 1 0 23760 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1867
timestamp 1626908933
transform 1 0 23856 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2349
timestamp 1626908933
transform 1 0 23760 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3802
timestamp 1626908933
transform 1 0 23856 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_142
timestamp 1626908933
transform 1 0 24384 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_740
timestamp 1626908933
transform 1 0 24384 0 -1 17316
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1800
timestamp 1626908933
transform 1 0 24048 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3735
timestamp 1626908933
transform 1 0 24048 0 1 16095
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_505
timestamp 1626908933
transform 1 0 24768 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1106
timestamp 1626908933
transform 1 0 24768 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1831
timestamp 1626908933
transform 1 0 24816 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3798
timestamp 1626908933
transform 1 0 24816 0 1 16539
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_83
timestamp 1626908933
transform 1 0 24500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_731
timestamp 1626908933
transform 1 0 24500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_83
timestamp 1626908933
transform 1 0 24500 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_731
timestamp 1626908933
transform 1 0 24500 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_13
timestamp 1626908933
transform 1 0 22560 0 -1 17316
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_1
timestamp 1626908933
transform 1 0 22560 0 -1 17316
box -38 -49 1862 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_862
timestamp 1626908933
transform 1 0 24960 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1853
timestamp 1626908933
transform 1 0 24960 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1800
timestamp 1626908933
transform 1 0 25872 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3767
timestamp 1626908933
transform 1 0 25872 0 1 16095
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1818
timestamp 1626908933
transform 1 0 25872 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3753
timestamp 1626908933
transform 1 0 25872 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_387
timestamp 1626908933
transform 1 0 25968 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2322
timestamp 1626908933
transform 1 0 25968 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_412
timestamp 1626908933
transform 1 0 26256 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2347
timestamp 1626908933
transform 1 0 26256 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_363
timestamp 1626908933
transform 1 0 26448 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1894
timestamp 1626908933
transform 1 0 26352 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2330
timestamp 1626908933
transform 1 0 26448 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3861
timestamp 1626908933
transform 1 0 26352 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1799
timestamp 1626908933
transform 1 0 26544 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1865
timestamp 1626908933
transform 1 0 26352 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3734
timestamp 1626908933
transform 1 0 26544 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3800
timestamp 1626908933
transform 1 0 26352 0 1 16317
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_707
timestamp 1626908933
transform 1 0 26900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_59
timestamp 1626908933
transform 1 0 26900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_707
timestamp 1626908933
transform 1 0 26900 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_59
timestamp 1626908933
transform 1 0 26900 0 1 16650
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3764
timestamp 1626908933
transform 1 0 26736 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1797
timestamp 1626908933
transform 1 0 26736 0 1 16095
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1307
timestamp 1626908933
transform 1 0 26880 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_316
timestamp 1626908933
transform 1 0 26880 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_689
timestamp 1626908933
transform 1 0 26976 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_91
timestamp 1626908933
transform 1 0 26976 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_169
timestamp 1626908933
transform 1 0 27456 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_526
timestamp 1626908933
transform 1 0 27456 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_77
timestamp 1626908933
transform 1 0 27648 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_675
timestamp 1626908933
transform 1 0 27648 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_314
timestamp 1626908933
transform 1 0 27552 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_315
timestamp 1626908933
transform 1 0 27360 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1305
timestamp 1626908933
transform 1 0 27552 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1306
timestamp 1626908933
transform 1 0 27360 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_14
timestamp 1626908933
transform -1 0 26880 0 -1 17316
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_2
timestamp 1626908933
transform -1 0 26880 0 -1 17316
box -38 -49 1862 715
use L1M1_PR  L1M1_PR_3362
timestamp 1626908933
transform 1 0 28176 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1427
timestamp 1626908933
transform 1 0 28176 0 1 16761
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3313
timestamp 1626908933
transform 1 0 28272 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1346
timestamp 1626908933
transform 1 0 28272 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_413
timestamp 1626908933
transform 1 0 29424 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2380
timestamp 1626908933
transform 1 0 29424 0 1 16243
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_35
timestamp 1626908933
transform 1 0 29300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_683
timestamp 1626908933
transform 1 0 29300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_35
timestamp 1626908933
transform 1 0 29300 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_683
timestamp 1626908933
transform 1 0 29300 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_162
timestamp 1626908933
transform 1 0 29856 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_763
timestamp 1626908933
transform 1 0 29856 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_313
timestamp 1626908933
transform 1 0 30048 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1304
timestamp 1626908933
transform 1 0 30048 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_45
timestamp 1626908933
transform 1 0 30144 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_767
timestamp 1626908933
transform 1 0 30144 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_15
timestamp 1626908933
transform -1 0 29856 0 -1 17316
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_3
timestamp 1626908933
transform -1 0 29856 0 -1 17316
box -38 -49 1862 715
use M1M2_PR  M1M2_PR_2374
timestamp 1626908933
transform 1 0 30864 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2373
timestamp 1626908933
transform 1 0 30864 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_407
timestamp 1626908933
transform 1 0 30864 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_406
timestamp 1626908933
transform 1 0 30864 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_0
timestamp 1626908933
transform 1 0 30912 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_69
timestamp 1626908933
transform 1 0 30912 0 -1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2337
timestamp 1626908933
transform 1 0 31056 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_402
timestamp 1626908933
transform 1 0 31056 0 1 16761
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1107
timestamp 1626908933
transform 1 0 31392 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_506
timestamp 1626908933
transform 1 0 31392 0 -1 17316
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_659
timestamp 1626908933
transform 1 0 31700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_11
timestamp 1626908933
transform 1 0 31700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_659
timestamp 1626908933
transform 1 0 31700 0 1 16650
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_11
timestamp 1626908933
transform 1 0 31700 0 1 16650
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1854
timestamp 1626908933
transform 1 0 31584 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_863
timestamp 1626908933
transform 1 0 31584 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1108
timestamp 1626908933
transform 1 0 31776 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_507
timestamp 1626908933
transform 1 0 31776 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_525
timestamp 1626908933
transform 1 0 31680 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_168
timestamp 1626908933
transform 1 0 31680 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_864
timestamp 1626908933
transform 1 0 31968 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1855
timestamp 1626908933
transform 1 0 31968 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1856
timestamp 1626908933
transform 1 0 192 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_865
timestamp 1626908933
transform 1 0 192 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1110
timestamp 1626908933
transform 1 0 384 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1109
timestamp 1626908933
transform 1 0 0 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_509
timestamp 1626908933
transform 1 0 384 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_508
timestamp 1626908933
transform 1 0 0 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_524
timestamp 1626908933
transform 1 0 288 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_167
timestamp 1626908933
transform 1 0 288 0 1 17316
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1283
timestamp 1626908933
transform 1 0 1700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_635
timestamp 1626908933
transform 1 0 1700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1283
timestamp 1626908933
transform 1 0 1700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_635
timestamp 1626908933
transform 1 0 1700 0 1 17316
box -100 -49 100 49
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_77
timestamp 1626908933
transform -1 0 3264 0 1 17316
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_31
timestamp 1626908933
transform -1 0 3264 0 1 17316
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1108
timestamp 1626908933
transform 1 0 3312 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3075
timestamp 1626908933
transform 1 0 3312 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1176
timestamp 1626908933
transform 1 0 3312 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3111
timestamp 1626908933
transform 1 0 3312 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1549
timestamp 1626908933
transform 1 0 3216 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3516
timestamp 1626908933
transform 1 0 3216 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1181
timestamp 1626908933
transform 1 0 3024 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1638
timestamp 1626908933
transform 1 0 3216 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3116
timestamp 1626908933
transform 1 0 3024 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3573
timestamp 1626908933
transform 1 0 3216 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1174
timestamp 1626908933
transform 1 0 3504 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3109
timestamp 1626908933
transform 1 0 3504 0 1 17057
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_611
timestamp 1626908933
transform 1 0 4100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1259
timestamp 1626908933
transform 1 0 4100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_611
timestamp 1626908933
transform 1 0 4100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1259
timestamp 1626908933
transform 1 0 4100 0 1 17316
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1548
timestamp 1626908933
transform 1 0 3216 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3515
timestamp 1626908933
transform 1 0 3216 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3110
timestamp 1626908933
transform 1 0 4368 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1175
timestamp 1626908933
transform 1 0 4368 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3108
timestamp 1626908933
transform 1 0 4560 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1173
timestamp 1626908933
transform 1 0 4560 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2368
timestamp 1626908933
transform 1 0 4656 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_401
timestamp 1626908933
transform 1 0 4656 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3881
timestamp 1626908933
transform 1 0 4368 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1914
timestamp 1626908933
transform 1 0 4368 0 1 17131
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3114
timestamp 1626908933
transform 1 0 4464 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1179
timestamp 1626908933
transform 1 0 4464 0 1 17205
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3078
timestamp 1626908933
transform 1 0 4560 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1111
timestamp 1626908933
transform 1 0 4560 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3170
timestamp 1626908933
transform 1 0 4368 0 1 17501
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1235
timestamp 1626908933
transform 1 0 4368 0 1 17501
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_166
timestamp 1626908933
transform 1 0 4992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_523
timestamp 1626908933
transform 1 0 4992 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1105
timestamp 1626908933
transform 1 0 4848 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3072
timestamp 1626908933
transform 1 0 4848 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_399
timestamp 1626908933
transform 1 0 5520 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1878
timestamp 1626908933
transform 1 0 5328 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2334
timestamp 1626908933
transform 1 0 5520 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3813
timestamp 1626908933
transform 1 0 5328 0 1 17131
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_603
timestamp 1626908933
transform 1 0 5088 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1325
timestamp 1626908933
transform 1 0 5088 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__a211oi_4  sky130_fd_sc_hs__a211oi_4_1
timestamp 1626908933
transform -1 0 4992 0 1 17316
box -38 -49 1766 715
use sky130_fd_sc_hs__a211oi_4  sky130_fd_sc_hs__a211oi_4_0
timestamp 1626908933
transform -1 0 4992 0 1 17316
box -38 -49 1766 715
use M1M2_PR  M1M2_PR_400
timestamp 1626908933
transform 1 0 5808 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2367
timestamp 1626908933
transform 1 0 5808 0 1 16909
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_55
timestamp 1626908933
transform 1 0 5856 0 1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_117
timestamp 1626908933
transform 1 0 5856 0 1 17316
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3789
timestamp 1626908933
transform 1 0 6384 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3785
timestamp 1626908933
transform 1 0 6288 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1854
timestamp 1626908933
transform 1 0 6384 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1850
timestamp 1626908933
transform 1 0 6288 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3841
timestamp 1626908933
transform 1 0 6288 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1874
timestamp 1626908933
transform 1 0 6288 0 1 16983
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1235
timestamp 1626908933
transform 1 0 6500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_587
timestamp 1626908933
transform 1 0 6500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1235
timestamp 1626908933
transform 1 0 6500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_587
timestamp 1626908933
transform 1 0 6500 0 1 17316
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3843
timestamp 1626908933
transform 1 0 6192 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1876
timestamp 1626908933
transform 1 0 6192 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_88
timestamp 1626908933
transform 1 0 6144 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_36
timestamp 1626908933
transform 1 0 6144 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_510
timestamp 1626908933
transform 1 0 6528 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1111
timestamp 1626908933
transform 1 0 6528 0 1 17316
box -38 -49 230 715
use L1M1_PR  L1M1_PR_466
timestamp 1626908933
transform 1 0 6576 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2401
timestamp 1626908933
transform 1 0 6576 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3788
timestamp 1626908933
transform 1 0 6672 0 1 17501
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1853
timestamp 1626908933
transform 1 0 6672 0 1 17501
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3846
timestamp 1626908933
transform 1 0 6672 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3845
timestamp 1626908933
transform 1 0 6672 0 1 17501
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1879
timestamp 1626908933
transform 1 0 6672 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1878
timestamp 1626908933
transform 1 0 6672 0 1 17501
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1857
timestamp 1626908933
transform 1 0 6720 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_866
timestamp 1626908933
transform 1 0 6720 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3784
timestamp 1626908933
transform 1 0 7056 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1849
timestamp 1626908933
transform 1 0 7056 0 1 17057
box -29 -23 29 23
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_43
timestamp 1626908933
transform 1 0 6816 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_18
timestamp 1626908933
transform 1 0 6816 0 1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3787
timestamp 1626908933
transform 1 0 7248 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2427
timestamp 1626908933
transform 1 0 7344 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1852
timestamp 1626908933
transform 1 0 7248 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_492
timestamp 1626908933
transform 1 0 7344 0 1 17131
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2466
timestamp 1626908933
transform 1 0 7344 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2465
timestamp 1626908933
transform 1 0 7344 0 1 17501
box -32 -32 32 32
use M1M2_PR  M1M2_PR_499
timestamp 1626908933
transform 1 0 7344 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_498
timestamp 1626908933
transform 1 0 7344 0 1 17501
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1112
timestamp 1626908933
transform 1 0 7680 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_511
timestamp 1626908933
transform 1 0 7680 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_89
timestamp 1626908933
transform 1 0 7296 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_37
timestamp 1626908933
transform 1 0 7296 0 1 17316
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3169
timestamp 1626908933
transform 1 0 7920 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1234
timestamp 1626908933
transform 1 0 7920 0 1 17427
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2434
timestamp 1626908933
transform 1 0 7920 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_467
timestamp 1626908933
transform 1 0 7920 0 1 17205
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1858
timestamp 1626908933
transform 1 0 7872 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_867
timestamp 1626908933
transform 1 0 7872 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__clkbuf_8  sky130_fd_sc_hs__clkbuf_8_0
timestamp 1626908933
transform 1 0 7968 0 1 17316
box -38 -49 1094 715
use sky130_fd_sc_hs__clkbuf_8  sky130_fd_sc_hs__clkbuf_8_1
timestamp 1626908933
transform 1 0 7968 0 1 17316
box -38 -49 1094 715
use M1M2_PR  M1M2_PR_3070
timestamp 1626908933
transform 1 0 8400 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1103
timestamp 1626908933
transform 1 0 8400 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3105
timestamp 1626908933
transform 1 0 8496 0 1 16835
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1170
timestamp 1626908933
transform 1 0 8496 0 1 16835
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2247
timestamp 1626908933
transform 1 0 8496 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_280
timestamp 1626908933
transform 1 0 8496 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3107
timestamp 1626908933
transform 1 0 8304 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1172
timestamp 1626908933
transform 1 0 8304 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2236
timestamp 1626908933
transform 1 0 8592 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_301
timestamp 1626908933
transform 1 0 8592 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3698
timestamp 1626908933
transform 1 0 8688 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1731
timestamp 1626908933
transform 1 0 8688 0 1 17427
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1211
timestamp 1626908933
transform 1 0 8900 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_563
timestamp 1626908933
transform 1 0 8900 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1211
timestamp 1626908933
transform 1 0 8900 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_563
timestamp 1626908933
transform 1 0 8900 0 1 17316
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3694
timestamp 1626908933
transform 1 0 8880 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3102
timestamp 1626908933
transform 1 0 8880 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1759
timestamp 1626908933
transform 1 0 8880 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1167
timestamp 1626908933
transform 1 0 8880 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3103
timestamp 1626908933
transform 1 0 9072 0 1 16835
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1168
timestamp 1626908933
transform 1 0 9072 0 1 16835
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3068
timestamp 1626908933
transform 1 0 9072 0 1 16835
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1101
timestamp 1626908933
transform 1 0 9072 0 1 16835
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1303
timestamp 1626908933
transform 1 0 9024 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_312
timestamp 1626908933
transform 1 0 9024 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_536
timestamp 1626908933
transform 1 0 9120 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1258
timestamp 1626908933
transform 1 0 9120 0 1 17316
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3100
timestamp 1626908933
transform 1 0 9552 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1165
timestamp 1626908933
transform 1 0 9552 0 1 17131
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3066
timestamp 1626908933
transform 1 0 9456 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1099
timestamp 1626908933
transform 1 0 9456 0 1 17131
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3098
timestamp 1626908933
transform 1 0 9264 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1163
timestamp 1626908933
transform 1 0 9264 0 1 17205
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3064
timestamp 1626908933
transform 1 0 9264 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1097
timestamp 1626908933
transform 1 0 9264 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2464
timestamp 1626908933
transform 1 0 9648 0 1 17501
box -32 -32 32 32
use M1M2_PR  M1M2_PR_497
timestamp 1626908933
transform 1 0 9648 0 1 17501
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_165
timestamp 1626908933
transform 1 0 9984 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_522
timestamp 1626908933
transform 1 0 9984 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_311
timestamp 1626908933
transform 1 0 9888 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1302
timestamp 1626908933
transform 1 0 9888 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_219
timestamp 1626908933
transform 1 0 10128 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_220
timestamp 1626908933
transform 1 0 10128 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2186
timestamp 1626908933
transform 1 0 10128 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2187
timestamp 1626908933
transform 1 0 10128 0 1 17205
box -32 -32 32 32
use sky130_fd_sc_hs__a222oi_1  sky130_fd_sc_hs__a222oi_1_0
timestamp 1626908933
transform 1 0 10080 0 1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__a222oi_1  sky130_fd_sc_hs__a222oi_1_2
timestamp 1626908933
transform 1 0 10080 0 1 17316
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1079
timestamp 1626908933
transform 1 0 10512 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3014
timestamp 1626908933
transform 1 0 10512 0 1 16909
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_310
timestamp 1626908933
transform 1 0 10944 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1301
timestamp 1626908933
transform 1 0 10944 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_275
timestamp 1626908933
transform 1 0 10800 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2242
timestamp 1626908933
transform 1 0 10800 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_237
timestamp 1626908933
transform 1 0 10704 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2172
timestamp 1626908933
transform 1 0 10704 0 1 17205
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_495
timestamp 1626908933
transform 1 0 11040 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1217
timestamp 1626908933
transform 1 0 11040 0 1 17316
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1082
timestamp 1626908933
transform 1 0 11280 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3017
timestamp 1626908933
transform 1 0 11280 0 1 17057
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_539
timestamp 1626908933
transform 1 0 11300 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1187
timestamp 1626908933
transform 1 0 11300 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_539
timestamp 1626908933
transform 1 0 11300 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1187
timestamp 1626908933
transform 1 0 11300 0 1 17316
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1010
timestamp 1626908933
transform 1 0 11664 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2977
timestamp 1626908933
transform 1 0 11664 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1075
timestamp 1626908933
transform 1 0 11664 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1078
timestamp 1626908933
transform 1 0 11472 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3010
timestamp 1626908933
transform 1 0 11664 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3013
timestamp 1626908933
transform 1 0 11472 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_309
timestamp 1626908933
transform 1 0 11808 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1300
timestamp 1626908933
transform 1 0 11808 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_51
timestamp 1626908933
transform -1 0 12192 0 1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_113
timestamp 1626908933
transform -1 0 12192 0 1 17316
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1012
timestamp 1626908933
transform 1 0 12144 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1016
timestamp 1626908933
transform 1 0 12048 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2979
timestamp 1626908933
transform 1 0 12144 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2983
timestamp 1626908933
transform 1 0 12048 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3586
timestamp 1626908933
transform 1 0 12528 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1619
timestamp 1626908933
transform 1 0 12528 0 1 17131
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2204
timestamp 1626908933
transform 1 0 12720 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2203
timestamp 1626908933
transform 1 0 12720 0 1 17501
box -29 -23 29 23
use L1M1_PR  L1M1_PR_269
timestamp 1626908933
transform 1 0 12720 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_268
timestamp 1626908933
transform 1 0 12720 0 1 17501
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2214
timestamp 1626908933
transform 1 0 12720 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2213
timestamp 1626908933
transform 1 0 12720 0 1 17501
box -32 -32 32 32
use M1M2_PR  M1M2_PR_247
timestamp 1626908933
transform 1 0 12720 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_246
timestamp 1626908933
transform 1 0 12720 0 1 17501
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1113
timestamp 1626908933
transform 1 0 12576 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_512
timestamp 1626908933
transform 1 0 12576 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_38
timestamp 1626908933
transform 1 0 12192 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_90
timestamp 1626908933
transform 1 0 12192 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_37
timestamp 1626908933
transform 1 0 13248 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_14
timestamp 1626908933
transform 1 0 13248 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_47
timestamp 1626908933
transform 1 0 12768 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_116
timestamp 1626908933
transform 1 0 12768 0 1 17316
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1163
timestamp 1626908933
transform 1 0 13700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_515
timestamp 1626908933
transform 1 0 13700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1163
timestamp 1626908933
transform 1 0 13700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_515
timestamp 1626908933
transform 1 0 13700 0 1 17316
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1054
timestamp 1626908933
transform 1 0 14064 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3021
timestamp 1626908933
transform 1 0 14064 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_161
timestamp 1626908933
transform 1 0 14400 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_762
timestamp 1626908933
transform 1 0 14400 0 1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1060
timestamp 1626908933
transform 1 0 14256 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3027
timestamp 1626908933
transform 1 0 14256 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1658
timestamp 1626908933
transform 1 0 14256 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3593
timestamp 1626908933
transform 1 0 14256 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_332
timestamp 1626908933
transform 1 0 14592 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_930
timestamp 1626908933
transform 1 0 14592 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_44
timestamp 1626908933
transform 1 0 14016 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_106
timestamp 1626908933
transform 1 0 14016 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_164
timestamp 1626908933
transform 1 0 14976 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_521
timestamp 1626908933
transform 1 0 14976 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1703
timestamp 1626908933
transform 1 0 14832 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3638
timestamp 1626908933
transform 1 0 14832 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3592
timestamp 1626908933
transform 1 0 15216 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1657
timestamp 1626908933
transform 1 0 15216 0 1 17057
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3536
timestamp 1626908933
transform 1 0 15216 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1569
timestamp 1626908933
transform 1 0 15216 0 1 17057
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3529
timestamp 1626908933
transform 1 0 15312 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1594
timestamp 1626908933
transform 1 0 15312 0 1 17057
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3474
timestamp 1626908933
transform 1 0 15408 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1507
timestamp 1626908933
transform 1 0 15408 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3631
timestamp 1626908933
transform 1 0 15120 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1664
timestamp 1626908933
transform 1 0 15120 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3535
timestamp 1626908933
transform 1 0 15216 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1568
timestamp 1626908933
transform 1 0 15216 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3473
timestamp 1626908933
transform 1 0 15408 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1506
timestamp 1626908933
transform 1 0 15408 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2904
timestamp 1626908933
transform 1 0 15504 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_937
timestamp 1626908933
transform 1 0 15504 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_319
timestamp 1626908933
transform 1 0 15072 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_917
timestamp 1626908933
transform 1 0 15072 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_31
timestamp 1626908933
transform 1 0 15456 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_93
timestamp 1626908933
transform 1 0 15456 0 1 17316
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1748
timestamp 1626908933
transform 1 0 15600 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3683
timestamp 1626908933
transform 1 0 15600 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1593
timestamp 1626908933
transform 1 0 15696 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3528
timestamp 1626908933
transform 1 0 15696 0 1 17427
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_491
timestamp 1626908933
transform 1 0 16100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1139
timestamp 1626908933
transform 1 0 16100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_491
timestamp 1626908933
transform 1 0 16100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1139
timestamp 1626908933
transform 1 0 16100 0 1 17316
box -100 -49 100 49
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_15
timestamp 1626908933
transform 1 0 15840 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_38
timestamp 1626908933
transform 1 0 15840 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1859
timestamp 1626908933
transform 1 0 16608 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_868
timestamp 1626908933
transform 1 0 16608 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3672
timestamp 1626908933
transform 1 0 16944 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2126
timestamp 1626908933
transform 1 0 16944 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1705
timestamp 1626908933
transform 1 0 16944 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_159
timestamp 1626908933
transform 1 0 16944 0 1 17427
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1299
timestamp 1626908933
transform 1 0 16992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_308
timestamp 1626908933
transform 1 0 16992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_95
timestamp 1626908933
transform -1 0 16992 0 1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_33
timestamp 1626908933
transform -1 0 16992 0 1 17316
box -38 -49 326 715
use M1M2_PR  M1M2_PR_940
timestamp 1626908933
transform 1 0 17040 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2907
timestamp 1626908933
transform 1 0 17040 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_368
timestamp 1626908933
transform 1 0 17088 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1090
timestamp 1626908933
transform 1 0 17088 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_28
timestamp 1626908933
transform 1 0 17856 0 1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_89
timestamp 1626908933
transform 1 0 17856 0 1 17316
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1456
timestamp 1626908933
transform 1 0 18192 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1661
timestamp 1626908933
transform 1 0 17904 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3423
timestamp 1626908933
transform 1 0 18192 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3628
timestamp 1626908933
transform 1 0 17904 0 1 17131
box -32 -32 32 32
use L1M1_PR  L1M1_PR_174
timestamp 1626908933
transform 1 0 18192 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1542
timestamp 1626908933
transform 1 0 17904 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2109
timestamp 1626908933
transform 1 0 18192 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3477
timestamp 1626908933
transform 1 0 17904 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_39
timestamp 1626908933
transform 1 0 18144 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_91
timestamp 1626908933
transform 1 0 18144 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_869
timestamp 1626908933
transform 1 0 18528 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1860
timestamp 1626908933
transform 1 0 18528 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1742
timestamp 1626908933
transform 1 0 18288 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3677
timestamp 1626908933
transform 1 0 18288 0 1 16983
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_467
timestamp 1626908933
transform 1 0 18500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1115
timestamp 1626908933
transform 1 0 18500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_467
timestamp 1626908933
transform 1 0 18500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1115
timestamp 1626908933
transform 1 0 18500 0 1 17316
box -100 -49 100 49
use M1M2_PR  M1M2_PR_756
timestamp 1626908933
transform 1 0 19056 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1702
timestamp 1626908933
transform 1 0 18768 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2723
timestamp 1626908933
transform 1 0 19056 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3669
timestamp 1626908933
transform 1 0 18768 0 1 16909
box -32 -32 32 32
use L1M1_PR  L1M1_PR_784
timestamp 1626908933
transform 1 0 18960 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2719
timestamp 1626908933
transform 1 0 18960 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_81
timestamp 1626908933
transform 1 0 18624 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_12
timestamp 1626908933
transform 1 0 18624 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_240
timestamp 1626908933
transform 1 0 19104 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_838
timestamp 1626908933
transform 1 0 19104 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_513
timestamp 1626908933
transform 1 0 19776 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1114
timestamp 1626908933
transform 1 0 19776 0 1 17316
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1008
timestamp 1626908933
transform 1 0 19632 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2943
timestamp 1626908933
transform 1 0 19632 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_32
timestamp 1626908933
transform -1 0 19776 0 1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_94
timestamp 1626908933
transform -1 0 19776 0 1 17316
box -38 -49 326 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_104
timestamp 1626908933
transform 1 0 20256 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_35
timestamp 1626908933
transform 1 0 20256 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_163
timestamp 1626908933
transform 1 0 19968 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_520
timestamp 1626908933
transform 1 0 19968 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_514
timestamp 1626908933
transform 1 0 20064 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1115
timestamp 1626908933
transform 1 0 20064 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_160
timestamp 1626908933
transform 1 0 20736 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_761
timestamp 1626908933
transform 1 0 20736 0 1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_367
timestamp 1626908933
transform 1 0 20496 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1692
timestamp 1626908933
transform 1 0 20592 0 1 16835
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2334
timestamp 1626908933
transform 1 0 20496 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3659
timestamp 1626908933
transform 1 0 20592 0 1 16835
box -32 -32 32 32
use M1M2_PR  M1M2_PR_163
timestamp 1626908933
transform 1 0 21456 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_946
timestamp 1626908933
transform 1 0 21072 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2130
timestamp 1626908933
transform 1 0 21456 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2913
timestamp 1626908933
transform 1 0 21072 0 1 17057
box -32 -32 32 32
use L1M1_PR  L1M1_PR_180
timestamp 1626908933
transform 1 0 21456 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1006
timestamp 1626908933
transform 1 0 21264 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2115
timestamp 1626908933
transform 1 0 21456 0 1 17057
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2941
timestamp 1626908933
transform 1 0 21264 0 1 17057
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1091
timestamp 1626908933
transform 1 0 20900 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_443
timestamp 1626908933
transform 1 0 20900 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1091
timestamp 1626908933
transform 1 0 20900 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_443
timestamp 1626908933
transform 1 0 20900 0 1 17316
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2912
timestamp 1626908933
transform 1 0 21072 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_945
timestamp 1626908933
transform 1 0 21072 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2129
timestamp 1626908933
transform 1 0 21456 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_162
timestamp 1626908933
transform 1 0 21456 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3622
timestamp 1626908933
transform 1 0 21648 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1655
timestamp 1626908933
transform 1 0 21648 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2113
timestamp 1626908933
transform 1 0 21744 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_178
timestamp 1626908933
transform 1 0 21744 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_282
timestamp 1626908933
transform 1 0 20928 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1004
timestamp 1626908933
transform 1 0 20928 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_40
timestamp 1626908933
transform -1 0 23904 0 1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_15
timestamp 1626908933
transform -1 0 23904 0 1 17316
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_2324
timestamp 1626908933
transform 1 0 22704 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_389
timestamp 1626908933
transform 1 0 22704 0 1 16909
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2331
timestamp 1626908933
transform 1 0 22992 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_364
timestamp 1626908933
transform 1 0 22992 0 1 16909
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1067
timestamp 1626908933
transform 1 0 23300 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_419
timestamp 1626908933
transform 1 0 23300 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1067
timestamp 1626908933
transform 1 0 23300 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_419
timestamp 1626908933
transform 1 0 23300 0 1 17316
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3296
timestamp 1626908933
transform 1 0 23376 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1361
timestamp 1626908933
transform 1 0 23376 0 1 16909
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3467
timestamp 1626908933
transform 1 0 23760 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1500
timestamp 1626908933
transform 1 0 23760 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_515
timestamp 1626908933
transform 1 0 23904 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1116
timestamp 1626908933
transform 1 0 23904 0 1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1272
timestamp 1626908933
transform 1 0 24048 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3239
timestamp 1626908933
transform 1 0 24048 0 1 16909
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1359
timestamp 1626908933
transform 1 0 24048 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3294
timestamp 1626908933
transform 1 0 24048 0 1 16909
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_870
timestamp 1626908933
transform 1 0 24096 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1861
timestamp 1626908933
transform 1 0 24096 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1342
timestamp 1626908933
transform 1 0 24240 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1343
timestamp 1626908933
transform 1 0 24240 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3309
timestamp 1626908933
transform 1 0 24240 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3310
timestamp 1626908933
transform 1 0 24240 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1424
timestamp 1626908933
transform 1 0 24240 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3359
timestamp 1626908933
transform 1 0 24240 0 1 17205
box -29 -23 29 23
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_7
timestamp 1626908933
transform 1 0 24192 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_32
timestamp 1626908933
transform 1 0 24192 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1862
timestamp 1626908933
transform 1 0 24864 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_871
timestamp 1626908933
transform 1 0 24864 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1117
timestamp 1626908933
transform 1 0 24672 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_516
timestamp 1626908933
transform 1 0 24672 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_519
timestamp 1626908933
transform 1 0 24960 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_162
timestamp 1626908933
transform 1 0 24960 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3361
timestamp 1626908933
transform 1 0 25200 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1426
timestamp 1626908933
transform 1 0 25200 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3295
timestamp 1626908933
transform 1 0 25392 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1360
timestamp 1626908933
transform 1 0 25392 0 1 16909
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3312
timestamp 1626908933
transform 1 0 25488 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3311
timestamp 1626908933
transform 1 0 25488 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1345
timestamp 1626908933
transform 1 0 25488 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1344
timestamp 1626908933
transform 1 0 25488 0 1 17427
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_395
timestamp 1626908933
transform 1 0 25700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1043
timestamp 1626908933
transform 1 0 25700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_395
timestamp 1626908933
transform 1 0 25700 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1043
timestamp 1626908933
transform 1 0 25700 0 1 17316
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1425
timestamp 1626908933
transform 1 0 25776 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3360
timestamp 1626908933
transform 1 0 25776 0 1 17427
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1423
timestamp 1626908933
transform 1 0 26064 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3390
timestamp 1626908933
transform 1 0 26064 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1804
timestamp 1626908933
transform 1 0 26256 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3771
timestamp 1626908933
transform 1 0 26256 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_34
timestamp 1626908933
transform 1 0 25824 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_9
timestamp 1626908933
transform 1 0 25824 0 1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_184
timestamp 1626908933
transform 1 0 25056 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_906
timestamp 1626908933
transform 1 0 25056 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_307
timestamp 1626908933
transform 1 0 26304 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1298
timestamp 1626908933
transform 1 0 26304 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_362
timestamp 1626908933
transform 1 0 26640 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2329
timestamp 1626908933
transform 1 0 26640 0 1 16909
box -32 -32 32 32
use L1M1_PR  L1M1_PR_386
timestamp 1626908933
transform 1 0 26736 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1363
timestamp 1626908933
transform 1 0 26448 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2321
timestamp 1626908933
transform 1 0 26736 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3298
timestamp 1626908933
transform 1 0 26448 0 1 16909
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_155
timestamp 1626908933
transform 1 0 26400 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_877
timestamp 1626908933
transform 1 0 26400 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_51
timestamp 1626908933
transform 1 0 27168 0 1 17316
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_5
timestamp 1626908933
transform 1 0 27168 0 1 17316
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1273
timestamp 1626908933
transform 1 0 28272 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3240
timestamp 1626908933
transform 1 0 28272 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1362
timestamp 1626908933
transform 1 0 28368 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3297
timestamp 1626908933
transform 1 0 28368 0 1 16909
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1297
timestamp 1626908933
transform 1 0 28464 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3264
timestamp 1626908933
transform 1 0 28464 0 1 17057
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_371
timestamp 1626908933
transform 1 0 28100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1019
timestamp 1626908933
transform 1 0 28100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_371
timestamp 1626908933
transform 1 0 28100 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1019
timestamp 1626908933
transform 1 0 28100 0 1 17316
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3299
timestamp 1626908933
transform 1 0 28656 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1364
timestamp 1626908933
transform 1 0 28656 0 1 16909
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_872
timestamp 1626908933
transform 1 0 29856 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1863
timestamp 1626908933
transform 1 0 29856 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_384
timestamp 1626908933
transform 1 0 29712 0 1 16909
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2319
timestamp 1626908933
transform 1 0 29712 0 1 16909
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_161
timestamp 1626908933
transform 1 0 29952 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_518
timestamp 1626908933
transform 1 0 29952 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_159
timestamp 1626908933
transform 1 0 30048 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_760
timestamp 1626908933
transform 1 0 30048 0 1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_358
timestamp 1626908933
transform 1 0 29904 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2325
timestamp 1626908933
transform 1 0 29904 0 1 16909
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1297
timestamp 1626908933
transform 1 0 30240 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_306
timestamp 1626908933
transform 1 0 30240 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_766
timestamp 1626908933
transform 1 0 30336 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_44
timestamp 1626908933
transform 1 0 30336 0 1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1884
timestamp 1626908933
transform 1 0 30672 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3851
timestamp 1626908933
transform 1 0 30672 0 1 16983
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_347
timestamp 1626908933
transform 1 0 30500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_995
timestamp 1626908933
transform 1 0 30500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_347
timestamp 1626908933
transform 1 0 30500 0 1 17316
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_995
timestamp 1626908933
transform 1 0 30500 0 1 17316
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_305
timestamp 1626908933
transform 1 0 31104 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1296
timestamp 1626908933
transform 1 0 31104 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_405
timestamp 1626908933
transform 1 0 30960 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2372
timestamp 1626908933
transform 1 0 30960 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_401
timestamp 1626908933
transform 1 0 31056 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1855
timestamp 1626908933
transform 1 0 30960 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2336
timestamp 1626908933
transform 1 0 31056 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3790
timestamp 1626908933
transform 1 0 30960 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_10
timestamp 1626908933
transform 1 0 31200 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_732
timestamp 1626908933
transform 1 0 31200 0 1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3769
timestamp 1626908933
transform 1 0 32016 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1802
timestamp 1626908933
transform 1 0 32016 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1864
timestamp 1626908933
transform 1 0 31968 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_873
timestamp 1626908933
transform 1 0 31968 0 1 17316
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_970
timestamp 1626908933
transform 1 0 500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_322
timestamp 1626908933
transform 1 0 500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_970
timestamp 1626908933
transform 1 0 500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_322
timestamp 1626908933
transform 1 0 500 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_759
timestamp 1626908933
transform 1 0 0 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_158
timestamp 1626908933
transform 1 0 0 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1432
timestamp 1626908933
transform 1 0 192 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_710
timestamp 1626908933
transform 1 0 192 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_304
timestamp 1626908933
transform 1 0 960 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1295
timestamp 1626908933
transform 1 0 960 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_286
timestamp 1626908933
transform 1 0 1008 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_287
timestamp 1626908933
transform 1 0 1008 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2253
timestamp 1626908933
transform 1 0 1008 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2254
timestamp 1626908933
transform 1 0 1008 0 1 17871
box -32 -32 32 32
use L1M1_PR  L1M1_PR_309
timestamp 1626908933
transform 1 0 1008 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2244
timestamp 1626908933
transform 1 0 1008 0 1 17871
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_676
timestamp 1626908933
transform 1 0 1440 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1398
timestamp 1626908933
transform 1 0 1440 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_572
timestamp 1626908933
transform 1 0 1056 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1170
timestamp 1626908933
transform 1 0 1056 0 -1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3142
timestamp 1626908933
transform 1 0 2064 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1175
timestamp 1626908933
transform 1 0 2064 0 1 17723
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1294
timestamp 1626908933
transform 1 0 2208 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_303
timestamp 1626908933
transform 1 0 2208 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1118
timestamp 1626908933
transform 1 0 2304 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_517
timestamp 1626908933
transform 1 0 2304 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_517
timestamp 1626908933
transform 1 0 2496 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_160
timestamp 1626908933
transform 1 0 2496 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3614
timestamp 1626908933
transform 1 0 2736 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1647
timestamp 1626908933
transform 1 0 2736 0 1 17649
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1119
timestamp 1626908933
transform 1 0 2592 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_518
timestamp 1626908933
transform 1 0 2592 0 -1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3662
timestamp 1626908933
transform 1 0 2832 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1727
timestamp 1626908933
transform 1 0 2832 0 1 17649
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_946
timestamp 1626908933
transform 1 0 2900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_298
timestamp 1626908933
transform 1 0 2900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_946
timestamp 1626908933
transform 1 0 2900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_298
timestamp 1626908933
transform 1 0 2900 0 1 17982
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2243
timestamp 1626908933
transform 1 0 2928 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_308
timestamp 1626908933
transform 1 0 2928 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3112
timestamp 1626908933
transform 1 0 3120 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1177
timestamp 1626908933
transform 1 0 3120 0 1 18093
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_302
timestamp 1626908933
transform 1 0 3264 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1293
timestamp 1626908933
transform 1 0 3264 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1107
timestamp 1626908933
transform 1 0 3312 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3074
timestamp 1626908933
transform 1 0 3312 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1236
timestamp 1626908933
transform 1 0 3504 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1637
timestamp 1626908933
transform 1 0 3216 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3171
timestamp 1626908933
transform 1 0 3504 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3572
timestamp 1626908933
transform 1 0 3216 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_121
timestamp 1626908933
transform -1 0 3264 0 -1 18648
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_52
timestamp 1626908933
transform -1 0 3264 0 -1 18648
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_645
timestamp 1626908933
transform 1 0 3360 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1367
timestamp 1626908933
transform 1 0 3360 0 -1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1179
timestamp 1626908933
transform 1 0 3696 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1913
timestamp 1626908933
transform 1 0 4368 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3146
timestamp 1626908933
transform 1 0 3696 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3880
timestamp 1626908933
transform 1 0 4368 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1240
timestamp 1626908933
transform 1 0 3696 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1881
timestamp 1626908933
transform 1 0 4080 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3175
timestamp 1626908933
transform 1 0 3696 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3816
timestamp 1626908933
transform 1 0 4080 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_305
timestamp 1626908933
transform 1 0 3888 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2272
timestamp 1626908933
transform 1 0 3888 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_328
timestamp 1626908933
transform 1 0 4272 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2263
timestamp 1626908933
transform 1 0 4272 0 1 18315
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_56
timestamp 1626908933
transform 1 0 4128 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_118
timestamp 1626908933
transform 1 0 4128 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_301
timestamp 1626908933
transform 1 0 4512 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1292
timestamp 1626908933
transform 1 0 4512 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_445
timestamp 1626908933
transform 1 0 4752 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_446
timestamp 1626908933
transform 1 0 4752 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2412
timestamp 1626908933
transform 1 0 4752 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2413
timestamp 1626908933
transform 1 0 4752 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_445
timestamp 1626908933
transform 1 0 4464 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2380
timestamp 1626908933
transform 1 0 4464 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1177
timestamp 1626908933
transform 1 0 4944 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3144
timestamp 1626908933
transform 1 0 4944 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1237
timestamp 1626908933
transform 1 0 4944 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3172
timestamp 1626908933
transform 1 0 4944 0 1 17649
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_274
timestamp 1626908933
transform 1 0 5300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_922
timestamp 1626908933
transform 1 0 5300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_274
timestamp 1626908933
transform 1 0 5300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_922
timestamp 1626908933
transform 1 0 5300 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_620
timestamp 1626908933
transform 1 0 4608 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1342
timestamp 1626908933
transform 1 0 4608 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_758
timestamp 1626908933
transform 1 0 5376 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_157
timestamp 1626908933
transform 1 0 5376 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_300
timestamp 1626908933
transform 1 0 5568 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1291
timestamp 1626908933
transform 1 0 5568 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_444
timestamp 1626908933
transform 1 0 5712 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_495
timestamp 1626908933
transform 1 0 5904 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1851
timestamp 1626908933
transform 1 0 5904 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2379
timestamp 1626908933
transform 1 0 5712 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2430
timestamp 1626908933
transform 1 0 5904 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3786
timestamp 1626908933
transform 1 0 5904 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2393
timestamp 1626908933
transform 1 0 6000 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_458
timestamp 1626908933
transform 1 0 6000 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2469
timestamp 1626908933
transform 1 0 6000 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_502
timestamp 1626908933
transform 1 0 6000 0 1 17797
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3764
timestamp 1626908933
transform 1 0 6000 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3204
timestamp 1626908933
transform 1 0 6288 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1829
timestamp 1626908933
transform 1 0 6000 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1269
timestamp 1626908933
transform 1 0 6288 0 1 18167
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3820
timestamp 1626908933
transform 1 0 6192 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1853
timestamp 1626908933
transform 1 0 6192 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_757
timestamp 1626908933
transform 1 0 6240 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_156
timestamp 1626908933
transform 1 0 6240 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_8
timestamp 1626908933
transform 1 0 5664 0 -1 18648
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_21
timestamp 1626908933
transform 1 0 5664 0 -1 18648
box -38 -49 614 715
use L1M1_PR  L1M1_PR_3783
timestamp 1626908933
transform 1 0 7056 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1848
timestamp 1626908933
transform 1 0 7056 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1290
timestamp 1626908933
transform 1 0 6432 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_299
timestamp 1626908933
transform 1 0 6432 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1297
timestamp 1626908933
transform 1 0 6528 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_575
timestamp 1626908933
transform 1 0 6528 0 -1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_457
timestamp 1626908933
transform 1 0 7344 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2424
timestamp 1626908933
transform 1 0 7344 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_482
timestamp 1626908933
transform 1 0 7344 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2417
timestamp 1626908933
transform 1 0 7344 0 1 17871
box -29 -23 29 23
use M1M2_PR  M1M2_PR_456
timestamp 1626908933
transform 1 0 7344 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2423
timestamp 1626908933
transform 1 0 7344 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_298
timestamp 1626908933
transform 1 0 7296 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_874
timestamp 1626908933
transform 1 0 7392 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1289
timestamp 1626908933
transform 1 0 7296 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1865
timestamp 1626908933
transform 1 0 7392 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_516
timestamp 1626908933
transform 1 0 7488 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_159
timestamp 1626908933
transform 1 0 7488 0 -1 18648
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_898
timestamp 1626908933
transform 1 0 7700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_250
timestamp 1626908933
transform 1 0 7700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_898
timestamp 1626908933
transform 1 0 7700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_250
timestamp 1626908933
transform 1 0 7700 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_155
timestamp 1626908933
transform 1 0 8064 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_756
timestamp 1626908933
transform 1 0 8064 0 -1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_303
timestamp 1626908933
transform 1 0 8016 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_457
timestamp 1626908933
transform 1 0 7824 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2238
timestamp 1626908933
transform 1 0 8016 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2392
timestamp 1626908933
transform 1 0 7824 0 1 18315
box -29 -23 29 23
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_1
timestamp 1626908933
transform 1 0 7584 0 -1 18648
box -38 -49 518 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_7
timestamp 1626908933
transform 1 0 7584 0 -1 18648
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1271
timestamp 1626908933
transform 1 0 8256 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_549
timestamp 1626908933
transform 1 0 8256 0 -1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_452
timestamp 1626908933
transform 1 0 8976 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2419
timestamp 1626908933
transform 1 0 8976 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_223
timestamp 1626908933
transform 1 0 9072 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_279
timestamp 1626908933
transform 1 0 8496 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2190
timestamp 1626908933
transform 1 0 9072 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2246
timestamp 1626908933
transform 1 0 8496 0 1 18241
box -32 -32 32 32
use L1M1_PR  L1M1_PR_243
timestamp 1626908933
transform 1 0 9072 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1268
timestamp 1626908933
transform 1 0 9072 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2178
timestamp 1626908933
transform 1 0 9072 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3203
timestamp 1626908933
transform 1 0 9072 0 1 18167
box -29 -23 29 23
use sky130_fd_sc_hs__a222oi_1  sky130_fd_sc_hs__a222oi_1_1
timestamp 1626908933
transform 1 0 9024 0 -1 18648
box -38 -49 902 715
use sky130_fd_sc_hs__a222oi_1  sky130_fd_sc_hs__a222oi_1_3
timestamp 1626908933
transform 1 0 9024 0 -1 18648
box -38 -49 902 715
use M1M2_PR  M1M2_PR_495
timestamp 1626908933
transform 1 0 9648 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_496
timestamp 1626908933
transform 1 0 9648 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2462
timestamp 1626908933
transform 1 0 9648 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2463
timestamp 1626908933
transform 1 0 9648 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_490
timestamp 1626908933
transform 1 0 9456 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2425
timestamp 1626908933
transform 1 0 9456 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2413
timestamp 1626908933
transform 1 0 9840 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_478
timestamp 1626908933
transform 1 0 9840 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2451
timestamp 1626908933
transform 1 0 9840 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2450
timestamp 1626908933
transform 1 0 9840 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_484
timestamp 1626908933
transform 1 0 9840 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_483
timestamp 1626908933
transform 1 0 9840 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_239
timestamp 1626908933
transform 1 0 10128 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_493
timestamp 1626908933
transform 1 0 10128 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2174
timestamp 1626908933
transform 1 0 10128 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2428
timestamp 1626908933
transform 1 0 10128 0 1 17797
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_226
timestamp 1626908933
transform 1 0 10100 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_874
timestamp 1626908933
transform 1 0 10100 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_226
timestamp 1626908933
transform 1 0 10100 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_874
timestamp 1626908933
transform 1 0 10100 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_297
timestamp 1626908933
transform 1 0 10080 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1288
timestamp 1626908933
transform 1 0 10080 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_755
timestamp 1626908933
transform 1 0 9888 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_154
timestamp 1626908933
transform 1 0 9888 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_513
timestamp 1626908933
transform 1 0 10176 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1235
timestamp 1626908933
transform 1 0 10176 0 -1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_491
timestamp 1626908933
transform 1 0 10416 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_492
timestamp 1626908933
transform 1 0 10416 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2458
timestamp 1626908933
transform 1 0 10416 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2459
timestamp 1626908933
transform 1 0 10416 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_451
timestamp 1626908933
transform 1 0 10320 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_487
timestamp 1626908933
transform 1 0 10512 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2386
timestamp 1626908933
transform 1 0 10320 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2422
timestamp 1626908933
transform 1 0 10512 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_241
timestamp 1626908933
transform 1 0 10896 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_270
timestamp 1626908933
transform 1 0 10608 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_297
timestamp 1626908933
transform 1 0 10800 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_477
timestamp 1626908933
transform 1 0 10896 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2176
timestamp 1626908933
transform 1 0 10896 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2205
timestamp 1626908933
transform 1 0 10608 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2232
timestamp 1626908933
transform 1 0 10800 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2412
timestamp 1626908933
transform 1 0 10896 0 1 17649
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_47
timestamp 1626908933
transform -1 0 11232 0 -1 18648
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_108
timestamp 1626908933
transform -1 0 11232 0 -1 18648
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_296
timestamp 1626908933
transform 1 0 11232 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1287
timestamp 1626908933
transform 1 0 11232 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_222
timestamp 1626908933
transform 1 0 11472 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2189
timestamp 1626908933
transform 1 0 11472 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1007
timestamp 1626908933
transform 1 0 11760 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2974
timestamp 1626908933
transform 1 0 11760 0 1 17649
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_482
timestamp 1626908933
transform 1 0 11712 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1204
timestamp 1626908933
transform 1 0 11712 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_393
timestamp 1626908933
transform 1 0 11328 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_991
timestamp 1626908933
transform 1 0 11328 0 -1 18648
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3008
timestamp 1626908933
transform 1 0 11952 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1073
timestamp 1626908933
transform 1 0 11952 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3012
timestamp 1626908933
transform 1 0 12144 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1077
timestamp 1626908933
transform 1 0 12144 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2978
timestamp 1626908933
transform 1 0 12144 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1011
timestamp 1626908933
transform 1 0 12144 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3016
timestamp 1626908933
transform 1 0 12048 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1081
timestamp 1626908933
transform 1 0 12048 0 1 17871
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2982
timestamp 1626908933
transform 1 0 12048 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1015
timestamp 1626908933
transform 1 0 12048 0 1 17871
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_158
timestamp 1626908933
transform 1 0 12480 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_515
timestamp 1626908933
transform 1 0 12480 0 -1 18648
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_202
timestamp 1626908933
transform 1 0 12500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_850
timestamp 1626908933
transform 1 0 12500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_202
timestamp 1626908933
transform 1 0 12500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_850
timestamp 1626908933
transform 1 0 12500 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_362
timestamp 1626908933
transform 1 0 12576 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_960
timestamp 1626908933
transform 1 0 12576 0 -1 18648
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3058
timestamp 1626908933
transform 1 0 13296 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1123
timestamp 1626908933
transform 1 0 13296 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3023
timestamp 1626908933
transform 1 0 13488 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1056
timestamp 1626908933
transform 1 0 13488 0 1 17649
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1183
timestamp 1626908933
transform 1 0 12960 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_461
timestamp 1626908933
transform 1 0 12960 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_754
timestamp 1626908933
transform 1 0 13728 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_153
timestamp 1626908933
transform 1 0 13728 0 -1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1119
timestamp 1626908933
transform 1 0 14064 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1121
timestamp 1626908933
transform 1 0 14160 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3054
timestamp 1626908933
transform 1 0 14064 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3056
timestamp 1626908933
transform 1 0 14160 0 1 17649
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_43
timestamp 1626908933
transform 1 0 14400 0 -1 18648
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_104
timestamp 1626908933
transform 1 0 14400 0 -1 18648
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_875
timestamp 1626908933
transform 1 0 14304 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1866
timestamp 1626908933
transform 1 0 14304 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1126
timestamp 1626908933
transform 1 0 14352 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3061
timestamp 1626908933
transform 1 0 14352 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_345
timestamp 1626908933
transform 1 0 13920 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_943
timestamp 1626908933
transform 1 0 13920 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_152
timestamp 1626908933
transform 1 0 14688 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_753
timestamp 1626908933
transform 1 0 14688 0 -1 18648
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_178
timestamp 1626908933
transform 1 0 14900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_826
timestamp 1626908933
transform 1 0 14900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_178
timestamp 1626908933
transform 1 0 14900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_826
timestamp 1626908933
transform 1 0 14900 0 1 17982
box -100 -49 100 49
use L1M1_PR  L1M1_PR_995
timestamp 1626908933
transform 1 0 15504 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2930
timestamp 1626908933
transform 1 0 15504 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_421
timestamp 1626908933
transform 1 0 14880 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1143
timestamp 1626908933
transform 1 0 14880 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_295
timestamp 1626908933
transform 1 0 15648 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1286
timestamp 1626908933
transform 1 0 15648 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_654
timestamp 1626908933
transform 1 0 15696 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2621
timestamp 1626908933
transform 1 0 15696 0 1 17723
box -32 -32 32 32
use L1M1_PR  L1M1_PR_668
timestamp 1626908933
transform 1 0 15600 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2603
timestamp 1626908933
transform 1 0 15600 0 1 17649
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_391
timestamp 1626908933
transform 1 0 16128 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1113
timestamp 1626908933
transform 1 0 16128 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_304
timestamp 1626908933
transform 1 0 15744 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_902
timestamp 1626908933
transform 1 0 15744 0 -1 18648
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2935
timestamp 1626908933
transform 1 0 16656 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2929
timestamp 1626908933
transform 1 0 16752 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2601
timestamp 1626908933
transform 1 0 16944 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1000
timestamp 1626908933
transform 1 0 16656 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_994
timestamp 1626908933
transform 1 0 16752 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_666
timestamp 1626908933
transform 1 0 16944 0 1 17649
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_154
timestamp 1626908933
transform 1 0 17300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_802
timestamp 1626908933
transform 1 0 17300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_154
timestamp 1626908933
transform 1 0 17300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_802
timestamp 1626908933
transform 1 0 17300 0 1 17982
box -100 -49 100 49
use M1M2_PR  M1M2_PR_939
timestamp 1626908933
transform 1 0 17040 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2906
timestamp 1626908933
transform 1 0 17040 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_999
timestamp 1626908933
transform 1 0 17040 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2934
timestamp 1626908933
transform 1 0 17040 0 1 18093
box -29 -23 29 23
use M1M2_PR  M1M2_PR_158
timestamp 1626908933
transform 1 0 16944 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2125
timestamp 1626908933
transform 1 0 16944 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_175
timestamp 1626908933
transform 1 0 16944 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2110
timestamp 1626908933
transform 1 0 16944 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1004
timestamp 1626908933
transform 1 0 17232 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2939
timestamp 1626908933
transform 1 0 17232 0 1 18315
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_57
timestamp 1626908933
transform -1 0 17472 0 -1 18648
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_18
timestamp 1626908933
transform -1 0 17472 0 -1 18648
box -38 -49 614 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_157
timestamp 1626908933
transform 1 0 17472 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_514
timestamp 1626908933
transform 1 0 17472 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_943
timestamp 1626908933
transform 1 0 17520 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_944
timestamp 1626908933
transform 1 0 17520 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2910
timestamp 1626908933
transform 1 0 17520 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2911
timestamp 1626908933
transform 1 0 17520 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1590
timestamp 1626908933
transform 1 0 17616 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3525
timestamp 1626908933
transform 1 0 17616 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_998
timestamp 1626908933
transform 1 0 17904 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2933
timestamp 1626908933
transform 1 0 17904 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2938
timestamp 1626908933
transform 1 0 18000 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1003
timestamp 1626908933
transform 1 0 18000 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3668
timestamp 1626908933
transform 1 0 18768 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2719
timestamp 1626908933
transform 1 0 19344 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1701
timestamp 1626908933
transform 1 0 18768 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_752
timestamp 1626908933
transform 1 0 19344 0 1 17797
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_39
timestamp 1626908933
transform 1 0 17568 0 -1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_14
timestamp 1626908933
transform 1 0 17568 0 -1 18648
box -38 -49 2246 715
use L1M1_PR  L1M1_PR_1002
timestamp 1626908933
transform 1 0 19536 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2937
timestamp 1626908933
transform 1 0 19536 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_161
timestamp 1626908933
transform 1 0 19920 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_942
timestamp 1626908933
transform 1 0 19824 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2128
timestamp 1626908933
transform 1 0 19920 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2909
timestamp 1626908933
transform 1 0 19824 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_780
timestamp 1626908933
transform 1 0 19824 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2715
timestamp 1626908933
transform 1 0 19824 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_176
timestamp 1626908933
transform 1 0 20304 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_778
timestamp 1626908933
transform 1 0 20400 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2111
timestamp 1626908933
transform 1 0 20304 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2713
timestamp 1626908933
transform 1 0 20400 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_177
timestamp 1626908933
transform 1 0 19728 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2112
timestamp 1626908933
transform 1 0 19728 0 1 18093
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_130
timestamp 1626908933
transform 1 0 19700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_778
timestamp 1626908933
transform 1 0 19700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_130
timestamp 1626908933
transform 1 0 19700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_778
timestamp 1626908933
transform 1 0 19700 0 1 17982
box -100 -49 100 49
use M1M2_PR  M1M2_PR_160
timestamp 1626908933
transform 1 0 19920 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2127
timestamp 1626908933
transform 1 0 19920 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1502
timestamp 1626908933
transform 1 0 20112 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3469
timestamp 1626908933
transform 1 0 20112 0 1 18241
box -32 -32 32 32
use L1M1_PR  L1M1_PR_390
timestamp 1626908933
transform 1 0 20208 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2325
timestamp 1626908933
transform 1 0 20208 0 1 18093
box -29 -23 29 23
use M1M2_PR  M1M2_PR_366
timestamp 1626908933
transform 1 0 20496 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2333
timestamp 1626908933
transform 1 0 20496 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1386
timestamp 1626908933
transform 1 0 21648 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3353
timestamp 1626908933
transform 1 0 21648 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1465
timestamp 1626908933
transform 1 0 22032 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3400
timestamp 1626908933
transform 1 0 22032 0 1 18315
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_106
timestamp 1626908933
transform 1 0 22100 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_754
timestamp 1626908933
transform 1 0 22100 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_106
timestamp 1626908933
transform 1 0 22100 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_754
timestamp 1626908933
transform 1 0 22100 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_62
timestamp 1626908933
transform -1 0 22464 0 -1 18648
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_16
timestamp 1626908933
transform -1 0 22464 0 -1 18648
box -38 -49 2726 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_156
timestamp 1626908933
transform 1 0 22464 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_513
timestamp 1626908933
transform 1 0 22464 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_390
timestamp 1626908933
transform 1 0 22128 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2357
timestamp 1626908933
transform 1 0 22128 0 1 18241
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1482
timestamp 1626908933
transform 1 0 22416 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3417
timestamp 1626908933
transform 1 0 22416 0 1 18241
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_151
timestamp 1626908933
transform 1 0 23328 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_752
timestamp 1626908933
transform 1 0 23328 0 -1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1689
timestamp 1626908933
transform 1 0 23088 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3656
timestamp 1626908933
transform 1 0 23088 0 1 17649
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_248
timestamp 1626908933
transform 1 0 22560 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_970
timestamp 1626908933
transform 1 0 22560 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_158
timestamp 1626908933
transform 1 0 23520 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_756
timestamp 1626908933
transform 1 0 23520 0 -1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1425
timestamp 1626908933
transform 1 0 23760 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3392
timestamp 1626908933
transform 1 0 23760 0 1 17723
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1587
timestamp 1626908933
transform 1 0 23856 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1738
timestamp 1626908933
transform 1 0 23568 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3522
timestamp 1626908933
transform 1 0 23856 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3673
timestamp 1626908933
transform 1 0 23568 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3358
timestamp 1626908933
transform 1 0 24240 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1423
timestamp 1626908933
transform 1 0 24240 0 1 17575
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3366
timestamp 1626908933
transform 1 0 24336 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3365
timestamp 1626908933
transform 1 0 24336 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1399
timestamp 1626908933
transform 1 0 24336 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1398
timestamp 1626908933
transform 1 0 24336 0 1 18241
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_730
timestamp 1626908933
transform 1 0 24500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_82
timestamp 1626908933
transform 1 0 24500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_730
timestamp 1626908933
transform 1 0 24500 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_82
timestamp 1626908933
transform 1 0 24500 0 1 17982
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3445
timestamp 1626908933
transform 1 0 24432 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1510
timestamp 1626908933
transform 1 0 24432 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3416
timestamp 1626908933
transform 1 0 24624 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1481
timestamp 1626908933
transform 1 0 24624 0 1 17871
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1867
timestamp 1626908933
transform 1 0 24672 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_876
timestamp 1626908933
transform 1 0 24672 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3419
timestamp 1626908933
transform 1 0 24816 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1484
timestamp 1626908933
transform 1 0 24816 0 1 18241
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_218
timestamp 1626908933
transform 1 0 23904 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_940
timestamp 1626908933
transform 1 0 23904 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_60
timestamp 1626908933
transform 1 0 24768 0 -1 18648
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_14
timestamp 1626908933
transform 1 0 24768 0 -1 18648
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3396
timestamp 1626908933
transform 1 0 25200 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1461
timestamp 1626908933
transform 1 0 25200 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3368
timestamp 1626908933
transform 1 0 24912 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3367
timestamp 1626908933
transform 1 0 24912 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3348
timestamp 1626908933
transform 1 0 25488 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1401
timestamp 1626908933
transform 1 0 24912 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1400
timestamp 1626908933
transform 1 0 24912 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1381
timestamp 1626908933
transform 1 0 25488 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3444
timestamp 1626908933
transform 1 0 26064 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3418
timestamp 1626908933
transform 1 0 26256 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1509
timestamp 1626908933
transform 1 0 26064 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1483
timestamp 1626908933
transform 1 0 26256 0 1 17871
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2352
timestamp 1626908933
transform 1 0 26544 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2351
timestamp 1626908933
transform 1 0 26544 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_385
timestamp 1626908933
transform 1 0 26544 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_384
timestamp 1626908933
transform 1 0 26544 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1405
timestamp 1626908933
transform 1 0 27312 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3372
timestamp 1626908933
transform 1 0 27312 0 1 17723
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1488
timestamp 1626908933
transform 1 0 27216 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3423
timestamp 1626908933
transform 1 0 27216 0 1 17723
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_58
timestamp 1626908933
transform 1 0 26900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_706
timestamp 1626908933
transform 1 0 26900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_58
timestamp 1626908933
transform 1 0 26900 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_706
timestamp 1626908933
transform 1 0 26900 0 1 17982
box -100 -49 100 49
use M1M2_PR  M1M2_PR_361
timestamp 1626908933
transform 1 0 26640 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2328
timestamp 1626908933
transform 1 0 26640 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_385
timestamp 1626908933
transform 1 0 27024 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2320
timestamp 1626908933
transform 1 0 27024 0 1 18093
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1404
timestamp 1626908933
transform 1 0 27312 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3371
timestamp 1626908933
transform 1 0 27312 0 1 18093
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1285
timestamp 1626908933
transform 1 0 27552 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_294
timestamp 1626908933
transform 1 0 27552 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_512
timestamp 1626908933
transform 1 0 27456 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_155
timestamp 1626908933
transform 1 0 27456 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3391
timestamp 1626908933
transform 1 0 27600 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1456
timestamp 1626908933
transform 1 0 27600 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3340
timestamp 1626908933
transform 1 0 27600 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3339
timestamp 1626908933
transform 1 0 27600 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1373
timestamp 1626908933
transform 1 0 27600 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1372
timestamp 1626908933
transform 1 0 27600 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_125
timestamp 1626908933
transform 1 0 27648 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_847
timestamp 1626908933
transform 1 0 27648 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_33
timestamp 1626908933
transform 1 0 28416 0 -1 18648
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_8
timestamp 1626908933
transform 1 0 28416 0 -1 18648
box -38 -49 518 715
use M1M2_PR  M1M2_PR_3773
timestamp 1626908933
transform 1 0 27792 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2343
timestamp 1626908933
transform 1 0 27888 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1806
timestamp 1626908933
transform 1 0 27792 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_376
timestamp 1626908933
transform 1 0 27888 0 1 17723
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_293
timestamp 1626908933
transform 1 0 28896 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1284
timestamp 1626908933
transform 1 0 28896 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1487
timestamp 1626908933
transform 1 0 28848 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3422
timestamp 1626908933
transform 1 0 28848 0 1 18093
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_34
timestamp 1626908933
transform 1 0 29300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_682
timestamp 1626908933
transform 1 0 29300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_34
timestamp 1626908933
transform 1 0 29300 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_682
timestamp 1626908933
transform 1 0 29300 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_90
timestamp 1626908933
transform 1 0 28992 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_812
timestamp 1626908933
transform 1 0 28992 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_20
timestamp 1626908933
transform 1 0 30144 0 -1 18648
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_5
timestamp 1626908933
transform 1 0 30144 0 -1 18648
box -38 -49 710 715
use L1M1_PR  L1M1_PR_2316
timestamp 1626908933
transform 1 0 29424 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_381
timestamp 1626908933
transform 1 0 29424 0 1 17871
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2322
timestamp 1626908933
transform 1 0 29520 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_355
timestamp 1626908933
transform 1 0 29520 0 1 17871
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_628
timestamp 1626908933
transform 1 0 29760 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_30
timestamp 1626908933
transform 1 0 29760 0 -1 18648
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3751
timestamp 1626908933
transform 1 0 30288 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1816
timestamp 1626908933
transform 1 0 30288 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3795
timestamp 1626908933
transform 1 0 30576 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2342
timestamp 1626908933
transform 1 0 30480 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1860
timestamp 1626908933
transform 1 0 30576 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_407
timestamp 1626908933
transform 1 0 30480 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3850
timestamp 1626908933
transform 1 0 30672 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1883
timestamp 1626908933
transform 1 0 30672 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3732
timestamp 1626908933
transform 1 0 30768 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1797
timestamp 1626908933
transform 1 0 30768 0 1 18093
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1283
timestamp 1626908933
transform 1 0 30816 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_292
timestamp 1626908933
transform 1 0 30816 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_404
timestamp 1626908933
transform 1 0 30960 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2371
timestamp 1626908933
transform 1 0 30960 0 1 18241
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_27
timestamp 1626908933
transform 1 0 30912 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_749
timestamp 1626908933
transform 1 0 30912 0 -1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1791
timestamp 1626908933
transform 1 0 31344 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3758
timestamp 1626908933
transform 1 0 31344 0 1 18093
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_154
timestamp 1626908933
transform 1 0 31680 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_511
timestamp 1626908933
transform 1 0 31680 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_519
timestamp 1626908933
transform 1 0 31776 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1120
timestamp 1626908933
transform 1 0 31776 0 -1 18648
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_10
timestamp 1626908933
transform 1 0 31700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_658
timestamp 1626908933
transform 1 0 31700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_10
timestamp 1626908933
transform 1 0 31700 0 1 17982
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_658
timestamp 1626908933
transform 1 0 31700 0 1 17982
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_877
timestamp 1626908933
transform 1 0 31968 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1868
timestamp 1626908933
transform 1 0 31968 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1805
timestamp 1626908933
transform 1 0 31920 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3772
timestamp 1626908933
transform 1 0 31920 0 1 17797
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_520
timestamp 1626908933
transform 1 0 0 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1121
timestamp 1626908933
transform 1 0 0 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_878
timestamp 1626908933
transform 1 0 192 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1869
timestamp 1626908933
transform 1 0 192 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_153
timestamp 1626908933
transform 1 0 288 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_510
timestamp 1626908933
transform 1 0 288 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_521
timestamp 1626908933
transform 1 0 384 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1122
timestamp 1626908933
transform 1 0 384 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_879
timestamp 1626908933
transform 1 0 576 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1870
timestamp 1626908933
transform 1 0 576 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_330
timestamp 1626908933
transform 1 0 1008 0 1 18759
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2265
timestamp 1626908933
transform 1 0 1008 0 1 18759
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1282
timestamp 1626908933
transform 1 0 1700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_634
timestamp 1626908933
transform 1 0 1700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1282
timestamp 1626908933
transform 1 0 1700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_634
timestamp 1626908933
transform 1 0 1700 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3613
timestamp 1626908933
transform 1 0 2736 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3141
timestamp 1626908933
transform 1 0 2064 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1646
timestamp 1626908933
transform 1 0 2736 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1174
timestamp 1626908933
transform 1 0 2064 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_53
timestamp 1626908933
transform -1 0 3360 0 1 18648
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_7
timestamp 1626908933
transform -1 0 3360 0 1 18648
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_307
timestamp 1626908933
transform 1 0 3312 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2242
timestamp 1626908933
transform 1 0 3312 0 1 18537
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1539
timestamp 1626908933
transform 1 0 3312 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3506
timestamp 1626908933
transform 1 0 3312 0 1 19055
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1625
timestamp 1626908933
transform 1 0 3312 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1726
timestamp 1626908933
transform 1 0 2928 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3560
timestamp 1626908933
transform 1 0 3312 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3661
timestamp 1626908933
transform 1 0 2928 0 1 18981
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_644
timestamp 1626908933
transform 1 0 3360 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1366
timestamp 1626908933
transform 1 0 3360 0 1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_306
timestamp 1626908933
transform 1 0 3792 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2273
timestamp 1626908933
transform 1 0 3792 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_474
timestamp 1626908933
transform 1 0 4176 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2441
timestamp 1626908933
transform 1 0 4176 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_470
timestamp 1626908933
transform 1 0 4176 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2405
timestamp 1626908933
transform 1 0 4176 0 1 18389
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_610
timestamp 1626908933
transform 1 0 4100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1258
timestamp 1626908933
transform 1 0 4100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_610
timestamp 1626908933
transform 1 0 4100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1258
timestamp 1626908933
transform 1 0 4100 0 1 18648
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_291
timestamp 1626908933
transform 1 0 4128 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1282
timestamp 1626908933
transform 1 0 4128 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3177
timestamp 1626908933
transform 1 0 4368 0 1 18463
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1242
timestamp 1626908933
transform 1 0 4368 0 1 18463
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3148
timestamp 1626908933
transform 1 0 4368 0 1 18463
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2440
timestamp 1626908933
transform 1 0 4272 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1181
timestamp 1626908933
transform 1 0 4368 0 1 18463
box -32 -32 32 32
use M1M2_PR  M1M2_PR_473
timestamp 1626908933
transform 1 0 4272 0 1 18759
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_619
timestamp 1626908933
transform 1 0 4224 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1341
timestamp 1626908933
transform 1 0 4224 0 1 18648
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3202
timestamp 1626908933
transform 1 0 4464 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1267
timestamp 1626908933
transform 1 0 4464 0 1 18389
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_751
timestamp 1626908933
transform 1 0 5088 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_150
timestamp 1626908933
transform 1 0 5088 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1324
timestamp 1626908933
transform 1 0 5280 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_602
timestamp 1626908933
transform 1 0 5280 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_509
timestamp 1626908933
transform 1 0 4992 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_152
timestamp 1626908933
transform 1 0 4992 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3201
timestamp 1626908933
transform 1 0 5808 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1266
timestamp 1626908933
transform 1 0 5808 0 1 18389
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2468
timestamp 1626908933
transform 1 0 6000 0 1 18463
box -32 -32 32 32
use M1M2_PR  M1M2_PR_501
timestamp 1626908933
transform 1 0 6000 0 1 18463
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1088
timestamp 1626908933
transform 1 0 6048 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_490
timestamp 1626908933
transform 1 0 6048 0 1 18648
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1234
timestamp 1626908933
transform 1 0 6500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_586
timestamp 1626908933
transform 1 0 6500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1234
timestamp 1626908933
transform 1 0 6500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_586
timestamp 1626908933
transform 1 0 6500 0 1 18648
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1281
timestamp 1626908933
transform 1 0 6432 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_290
timestamp 1626908933
transform 1 0 6432 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1296
timestamp 1626908933
transform 1 0 6528 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_574
timestamp 1626908933
transform 1 0 6528 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_149
timestamp 1626908933
transform 1 0 7296 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_750
timestamp 1626908933
transform 1 0 7296 0 1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_285
timestamp 1626908933
transform 1 0 7344 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1634
timestamp 1626908933
transform 1 0 7536 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2252
timestamp 1626908933
transform 1 0 7344 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3601
timestamp 1626908933
transform 1 0 7536 0 1 18981
box -32 -32 32 32
use L1M1_PR  L1M1_PR_465
timestamp 1626908933
transform 1 0 7632 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2400
timestamp 1626908933
transform 1 0 7632 0 1 18389
box -29 -23 29 23
use M1M2_PR  M1M2_PR_465
timestamp 1626908933
transform 1 0 7920 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_466
timestamp 1626908933
transform 1 0 7920 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2432
timestamp 1626908933
transform 1 0 7920 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2433
timestamp 1626908933
transform 1 0 7920 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_447
timestamp 1626908933
transform 1 0 8016 0 1 18463
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2382
timestamp 1626908933
transform 1 0 8016 0 1 18463
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_555
timestamp 1626908933
transform 1 0 7872 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1277
timestamp 1626908933
transform 1 0 7872 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_466
timestamp 1626908933
transform 1 0 7488 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1064
timestamp 1626908933
transform 1 0 7488 0 1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2415
timestamp 1626908933
transform 1 0 8112 0 1 18463
box -32 -32 32 32
use M1M2_PR  M1M2_PR_448
timestamp 1626908933
transform 1 0 8112 0 1 18463
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_289
timestamp 1626908933
transform 1 0 8640 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1280
timestamp 1626908933
transform 1 0 8640 0 1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_451
timestamp 1626908933
transform 1 0 8976 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_464
timestamp 1626908933
transform 1 0 9072 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2418
timestamp 1626908933
transform 1 0 8976 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2431
timestamp 1626908933
transform 1 0 9072 0 1 18981
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_562
timestamp 1626908933
transform 1 0 8900 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1210
timestamp 1626908933
transform 1 0 8900 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_562
timestamp 1626908933
transform 1 0 8900 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1210
timestamp 1626908933
transform 1 0 8900 0 1 18648
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_535
timestamp 1626908933
transform 1 0 9120 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1257
timestamp 1626908933
transform 1 0 9120 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_445
timestamp 1626908933
transform 1 0 8736 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1043
timestamp 1626908933
transform 1 0 8736 0 1 18648
box -38 -49 422 715
use L1M1_PR  L1M1_PR_454
timestamp 1626908933
transform 1 0 9264 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2389
timestamp 1626908933
transform 1 0 9264 0 1 18389
box -29 -23 29 23
use M1M2_PR  M1M2_PR_252
timestamp 1626908933
transform 1 0 9552 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2219
timestamp 1626908933
transform 1 0 9552 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_274
timestamp 1626908933
transform 1 0 9552 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2209
timestamp 1626908933
transform 1 0 9552 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_300
timestamp 1626908933
transform 1 0 9744 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2235
timestamp 1626908933
transform 1 0 9744 0 1 18389
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_151
timestamp 1626908933
transform 1 0 9984 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_508
timestamp 1626908933
transform 1 0 9984 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_880
timestamp 1626908933
transform 1 0 9888 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1871
timestamp 1626908933
transform 1 0 9888 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1019
timestamp 1626908933
transform 1 0 10080 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_421
timestamp 1626908933
transform 1 0 10080 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1234
timestamp 1626908933
transform 1 0 10464 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_512
timestamp 1626908933
transform 1 0 10464 0 1 18648
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3022
timestamp 1626908933
transform 1 0 10992 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1087
timestamp 1626908933
transform 1 0 10992 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1083
timestamp 1626908933
transform 1 0 11184 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3018
timestamp 1626908933
transform 1 0 11184 0 1 18389
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_538
timestamp 1626908933
transform 1 0 11300 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1186
timestamp 1626908933
transform 1 0 11300 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_538
timestamp 1626908933
transform 1 0 11300 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1186
timestamp 1626908933
transform 1 0 11300 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_221
timestamp 1626908933
transform 1 0 11472 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2188
timestamp 1626908933
transform 1 0 11472 0 1 18981
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_481
timestamp 1626908933
transform 1 0 11232 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1203
timestamp 1626908933
transform 1 0 11232 0 1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1014
timestamp 1626908933
transform 1 0 12048 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1018
timestamp 1626908933
transform 1 0 12528 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2981
timestamp 1626908933
transform 1 0 12048 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2985
timestamp 1626908933
transform 1 0 12528 0 1 18537
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2175
timestamp 1626908933
transform 1 0 12048 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_240
timestamp 1626908933
transform 1 0 12048 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3015
timestamp 1626908933
transform 1 0 12144 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1080
timestamp 1626908933
transform 1 0 12144 0 1 18981
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2980
timestamp 1626908933
transform 1 0 12144 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1013
timestamp 1626908933
transform 1 0 12144 0 1 18981
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3019
timestamp 1626908933
transform 1 0 12336 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1084
timestamp 1626908933
transform 1 0 12336 0 1 18981
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2984
timestamp 1626908933
transform 1 0 12528 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1017
timestamp 1626908933
transform 1 0 12528 0 1 18981
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_361
timestamp 1626908933
transform 1 0 12576 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_959
timestamp 1626908933
transform 1 0 12576 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_27
timestamp 1626908933
transform -1 0 12576 0 1 18648
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_66
timestamp 1626908933
transform -1 0 12576 0 1 18648
box -38 -49 614 715
use M1M2_PR  M1M2_PR_3776
timestamp 1626908933
transform 1 0 13200 0 1 18833
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3030
timestamp 1626908933
transform 1 0 13296 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1809
timestamp 1626908933
transform 1 0 13200 0 1 18833
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1063
timestamp 1626908933
transform 1 0 13296 0 1 18537
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1182
timestamp 1626908933
transform 1 0 12960 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_460
timestamp 1626908933
transform 1 0 12960 0 1 18648
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1162
timestamp 1626908933
transform 1 0 13700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_514
timestamp 1626908933
transform 1 0 13700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1162
timestamp 1626908933
transform 1 0 13700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_514
timestamp 1626908933
transform 1 0 13700 0 1 18648
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1279
timestamp 1626908933
transform 1 0 13728 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_288
timestamp 1626908933
transform 1 0 13728 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_942
timestamp 1626908933
transform 1 0 13824 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_344
timestamp 1626908933
transform 1 0 13824 0 1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3026
timestamp 1626908933
transform 1 0 14256 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1059
timestamp 1626908933
transform 1 0 14256 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3060
timestamp 1626908933
transform 1 0 14448 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1125
timestamp 1626908933
transform 1 0 14448 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2208
timestamp 1626908933
transform 1 0 14640 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_273
timestamp 1626908933
transform 1 0 14640 0 1 18389
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2217
timestamp 1626908933
transform 1 0 14640 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_250
timestamp 1626908933
transform 1 0 14640 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3064
timestamp 1626908933
transform 1 0 14640 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1129
timestamp 1626908933
transform 1 0 14640 0 1 18537
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1057
timestamp 1626908933
transform 1 0 14352 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3024
timestamp 1626908933
transform 1 0 14352 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_429
timestamp 1626908933
transform 1 0 14208 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1151
timestamp 1626908933
transform 1 0 14208 0 1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2215
timestamp 1626908933
transform 1 0 14832 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_248
timestamp 1626908933
transform 1 0 14832 0 1 18981
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1130
timestamp 1626908933
transform 1 0 15072 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_408
timestamp 1626908933
transform 1 0 15072 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_507
timestamp 1626908933
transform 1 0 14976 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_150
timestamp 1626908933
transform 1 0 14976 0 1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1062
timestamp 1626908933
transform 1 0 16272 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3029
timestamp 1626908933
transform 1 0 16272 0 1 18537
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_490
timestamp 1626908933
transform 1 0 16100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1138
timestamp 1626908933
transform 1 0 16100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_490
timestamp 1626908933
transform 1 0 16100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1138
timestamp 1626908933
transform 1 0 16100 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1061
timestamp 1626908933
transform 1 0 16272 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3028
timestamp 1626908933
transform 1 0 16272 0 1 18981
box -32 -32 32 32
use L1M1_PR  L1M1_PR_271
timestamp 1626908933
transform 1 0 15888 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1124
timestamp 1626908933
transform 1 0 15984 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1128
timestamp 1626908933
transform 1 0 16176 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2206
timestamp 1626908933
transform 1 0 15888 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3059
timestamp 1626908933
transform 1 0 15984 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3063
timestamp 1626908933
transform 1 0 16176 0 1 18981
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_31
timestamp 1626908933
transform -1 0 16416 0 1 18648
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_70
timestamp 1626908933
transform -1 0 16416 0 1 18648
box -38 -49 614 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_894
timestamp 1626908933
transform 1 0 16416 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_296
timestamp 1626908933
transform 1 0 16416 0 1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1505
timestamp 1626908933
transform 1 0 17424 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1660
timestamp 1626908933
transform 1 0 17904 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3472
timestamp 1626908933
transform 1 0 17424 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3627
timestamp 1626908933
transform 1 0 17904 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1592
timestamp 1626908933
transform 1 0 17424 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1744
timestamp 1626908933
transform 1 0 17904 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3527
timestamp 1626908933
transform 1 0 17424 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3679
timestamp 1626908933
transform 1 0 17904 0 1 18389
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2124
timestamp 1626908933
transform 1 0 16944 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_157
timestamp 1626908933
transform 1 0 16944 0 1 19055
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3526
timestamp 1626908933
transform 1 0 17520 0 1 18759
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1591
timestamp 1626908933
transform 1 0 17520 0 1 18759
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3471
timestamp 1626908933
transform 1 0 17424 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1504
timestamp 1626908933
transform 1 0 17424 0 1 18759
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3678
timestamp 1626908933
transform 1 0 17904 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1743
timestamp 1626908933
transform 1 0 17904 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3626
timestamp 1626908933
transform 1 0 17904 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1659
timestamp 1626908933
transform 1 0 17904 0 1 18907
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_379
timestamp 1626908933
transform 1 0 16800 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1101
timestamp 1626908933
transform 1 0 16800 0 1 18648
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1114
timestamp 1626908933
transform 1 0 18500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_466
timestamp 1626908933
transform 1 0 18500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1114
timestamp 1626908933
transform 1 0 18500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_466
timestamp 1626908933
transform 1 0 18500 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3667
timestamp 1626908933
transform 1 0 18768 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1700
timestamp 1626908933
transform 1 0 18768 0 1 18981
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_38
timestamp 1626908933
transform 1 0 17568 0 1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtn_1  sky130_fd_sc_hs__dfrtn_1_13
timestamp 1626908933
transform 1 0 17568 0 1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_522
timestamp 1626908933
transform 1 0 19776 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1123
timestamp 1626908933
transform 1 0 19776 0 1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_173
timestamp 1626908933
transform 1 0 19728 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2108
timestamp 1626908933
transform 1 0 19728 0 1 19055
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_149
timestamp 1626908933
transform 1 0 19968 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_506
timestamp 1626908933
transform 1 0 19968 0 1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_422
timestamp 1626908933
transform 1 0 20304 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1534
timestamp 1626908933
transform 1 0 20400 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2389
timestamp 1626908933
transform 1 0 20304 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3501
timestamp 1626908933
transform 1 0 20400 0 1 18907
box -32 -32 32 32
use L1M1_PR  L1M1_PR_419
timestamp 1626908933
transform 1 0 20208 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1621
timestamp 1626908933
transform 1 0 20400 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2354
timestamp 1626908933
transform 1 0 20208 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3556
timestamp 1626908933
transform 1 0 20400 0 1 18907
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1090
timestamp 1626908933
transform 1 0 20900 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_442
timestamp 1626908933
transform 1 0 20900 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1090
timestamp 1626908933
transform 1 0 20900 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_442
timestamp 1626908933
transform 1 0 20900 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2359
timestamp 1626908933
transform 1 0 21264 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_392
timestamp 1626908933
transform 1 0 21264 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_6
timestamp 1626908933
transform 1 0 20064 0 1 18648
box -38 -49 2438 715
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_2
timestamp 1626908933
transform 1 0 20064 0 1 18648
box -38 -49 2438 715
use M1M2_PR  M1M2_PR_2356
timestamp 1626908933
transform 1 0 22128 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_389
timestamp 1626908933
transform 1 0 22128 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1278
timestamp 1626908933
transform 1 0 22464 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_287
timestamp 1626908933
transform 1 0 22464 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_969
timestamp 1626908933
transform 1 0 22560 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_247
timestamp 1626908933
transform 1 0 22560 0 1 18648
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1066
timestamp 1626908933
transform 1 0 23300 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_418
timestamp 1626908933
transform 1 0 23300 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1066
timestamp 1626908933
transform 1 0 23300 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_418
timestamp 1626908933
transform 1 0 23300 0 1 18648
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_749
timestamp 1626908933
transform 1 0 23328 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_148
timestamp 1626908933
transform 1 0 23328 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_755
timestamp 1626908933
transform 1 0 23520 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_157
timestamp 1626908933
transform 1 0 23520 0 1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3364
timestamp 1626908933
transform 1 0 24240 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1397
timestamp 1626908933
transform 1 0 24240 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_939
timestamp 1626908933
transform 1 0 23904 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_217
timestamp 1626908933
transform 1 0 23904 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1277
timestamp 1626908933
transform 1 0 24672 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_286
timestamp 1626908933
transform 1 0 24672 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1124
timestamp 1626908933
transform 1 0 24768 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_523
timestamp 1626908933
transform 1 0 24768 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_148
timestamp 1626908933
transform 1 0 24960 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_505
timestamp 1626908933
transform 1 0 24960 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1479
timestamp 1626908933
transform 1 0 25104 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3414
timestamp 1626908933
transform 1 0 25104 0 1 19055
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1380
timestamp 1626908933
transform 1 0 25488 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3347
timestamp 1626908933
transform 1 0 25488 0 1 18981
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1459
timestamp 1626908933
transform 1 0 25488 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3394
timestamp 1626908933
transform 1 0 25488 0 1 18981
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_394
timestamp 1626908933
transform 1 0 25700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1042
timestamp 1626908933
transform 1 0 25700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_394
timestamp 1626908933
transform 1 0 25700 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1042
timestamp 1626908933
transform 1 0 25700 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1422
timestamp 1626908933
transform 1 0 26064 0 1 18463
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3389
timestamp 1626908933
transform 1 0 26064 0 1 18463
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2350
timestamp 1626908933
transform 1 0 26544 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_383
timestamp 1626908933
transform 1 0 26544 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_57
timestamp 1626908933
transform 1 0 25056 0 1 18648
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_11
timestamp 1626908933
transform 1 0 25056 0 1 18648
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1349
timestamp 1626908933
transform 1 0 28464 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3316
timestamp 1626908933
transform 1 0 28464 0 1 18389
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1429
timestamp 1626908933
transform 1 0 28464 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3364
timestamp 1626908933
transform 1 0 28464 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1504
timestamp 1626908933
transform 1 0 28656 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3439
timestamp 1626908933
transform 1 0 28656 0 1 18389
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_370
timestamp 1626908933
transform 1 0 28100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1018
timestamp 1626908933
transform 1 0 28100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_370
timestamp 1626908933
transform 1 0 28100 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1018
timestamp 1626908933
transform 1 0 28100 0 1 18648
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1348
timestamp 1626908933
transform 1 0 28464 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3315
timestamp 1626908933
transform 1 0 28464 0 1 18759
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1430
timestamp 1626908933
transform 1 0 27888 0 1 18759
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3365
timestamp 1626908933
transform 1 0 27888 0 1 18759
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1274
timestamp 1626908933
transform 1 0 28176 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3241
timestamp 1626908933
transform 1 0 28176 0 1 19055
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1365
timestamp 1626908933
transform 1 0 28080 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3300
timestamp 1626908933
transform 1 0 28080 0 1 19055
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1296
timestamp 1626908933
transform 1 0 28464 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3263
timestamp 1626908933
transform 1 0 28464 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1276
timestamp 1626908933
transform 1 0 28944 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3243
timestamp 1626908933
transform 1 0 28944 0 1 19055
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1367
timestamp 1626908933
transform 1 0 28944 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3302
timestamp 1626908933
transform 1 0 28944 0 1 19055
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_42
timestamp 1626908933
transform 1 0 29568 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_640
timestamp 1626908933
transform 1 0 29568 0 1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_356
timestamp 1626908933
transform 1 0 29424 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_357
timestamp 1626908933
transform 1 0 29424 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2323
timestamp 1626908933
transform 1 0 29424 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2324
timestamp 1626908933
transform 1 0 29424 0 1 18537
box -32 -32 32 32
use L1M1_PR  L1M1_PR_380
timestamp 1626908933
transform 1 0 29424 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2315
timestamp 1626908933
transform 1 0 29424 0 1 19055
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_147
timestamp 1626908933
transform 1 0 29952 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_504
timestamp 1626908933
transform 1 0 29952 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_147
timestamp 1626908933
transform 1 0 30048 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_748
timestamp 1626908933
transform 1 0 30048 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_285
timestamp 1626908933
transform 1 0 30240 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1276
timestamp 1626908933
transform 1 0 30240 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_379
timestamp 1626908933
transform 1 0 30192 0 1 18537
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2314
timestamp 1626908933
transform 1 0 30192 0 1 18537
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_43
timestamp 1626908933
transform 1 0 30336 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_765
timestamp 1626908933
transform 1 0 30336 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_16
timestamp 1626908933
transform -1 0 29568 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_4
timestamp 1626908933
transform -1 0 29568 0 1 18648
box -38 -49 1862 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_994
timestamp 1626908933
transform 1 0 30500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_346
timestamp 1626908933
transform 1 0 30500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_994
timestamp 1626908933
transform 1 0 30500 0 1 18648
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_346
timestamp 1626908933
transform 1 0 30500 0 1 18648
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1275
timestamp 1626908933
transform 1 0 31104 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_284
timestamp 1626908933
transform 1 0 31104 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_731
timestamp 1626908933
transform 1 0 31200 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_9
timestamp 1626908933
transform 1 0 31200 0 1 18648
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3794
timestamp 1626908933
transform 1 0 31536 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3775
timestamp 1626908933
transform 1 0 32016 0 1 18833
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1827
timestamp 1626908933
transform 1 0 31536 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1808
timestamp 1626908933
transform 1 0 32016 0 1 18833
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1872
timestamp 1626908933
transform 1 0 31968 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_881
timestamp 1626908933
transform 1 0 31968 0 1 18648
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_969
timestamp 1626908933
transform 1 0 500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_321
timestamp 1626908933
transform 1 0 500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_969
timestamp 1626908933
transform 1 0 500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_321
timestamp 1626908933
transform 1 0 500 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_747
timestamp 1626908933
transform 1 0 0 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_146
timestamp 1626908933
transform 1 0 0 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1431
timestamp 1626908933
transform 1 0 192 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_709
timestamp 1626908933
transform 1 0 192 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1274
timestamp 1626908933
transform 1 0 960 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_283
timestamp 1626908933
transform 1 0 960 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1169
timestamp 1626908933
transform 1 0 1056 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_571
timestamp 1626908933
transform 1 0 1056 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1397
timestamp 1626908933
transform 1 0 1440 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_675
timestamp 1626908933
transform 1 0 1440 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1273
timestamp 1626908933
transform 1 0 2208 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_282
timestamp 1626908933
transform 1 0 2208 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1125
timestamp 1626908933
transform 1 0 2304 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_524
timestamp 1626908933
transform 1 0 2304 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_503
timestamp 1626908933
transform 1 0 2496 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_146
timestamp 1626908933
transform 1 0 2496 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_10
timestamp 1626908933
transform 1 0 2688 0 -1 19980
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_2
timestamp 1626908933
transform 1 0 2688 0 -1 19980
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1873
timestamp 1626908933
transform 1 0 2592 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_882
timestamp 1626908933
transform 1 0 2592 0 -1 19980
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_945
timestamp 1626908933
transform 1 0 2900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_297
timestamp 1626908933
transform 1 0 2900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_945
timestamp 1626908933
transform 1 0 2900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_297
timestamp 1626908933
transform 1 0 2900 0 1 19314
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3561
timestamp 1626908933
transform 1 0 3120 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1626
timestamp 1626908933
transform 1 0 3120 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2977
timestamp 1626908933
transform 1 0 3024 0 1 19573
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2264
timestamp 1626908933
transform 1 0 3024 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1042
timestamp 1626908933
transform 1 0 3024 0 1 19573
box -29 -23 29 23
use L1M1_PR  L1M1_PR_329
timestamp 1626908933
transform 1 0 3024 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2946
timestamp 1626908933
transform 1 0 3120 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_979
timestamp 1626908933
transform 1 0 3120 0 1 19573
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_281
timestamp 1626908933
transform 1 0 3360 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1272
timestamp 1626908933
transform 1 0 3360 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1538
timestamp 1626908933
transform 1 0 3312 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3505
timestamp 1626908933
transform 1 0 3312 0 1 19425
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_535
timestamp 1626908933
transform 1 0 3456 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1133
timestamp 1626908933
transform 1 0 3456 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_280
timestamp 1626908933
transform 1 0 3840 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_883
timestamp 1626908933
transform 1 0 3936 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1271
timestamp 1626908933
transform 1 0 3840 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1874
timestamp 1626908933
transform 1 0 3936 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_304
timestamp 1626908933
transform 1 0 3888 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1178
timestamp 1626908933
transform 1 0 3696 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2271
timestamp 1626908933
transform 1 0 3888 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3145
timestamp 1626908933
transform 1 0 3696 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1180
timestamp 1626908933
transform 1 0 4368 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3147
timestamp 1626908933
transform 1 0 4368 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_446
timestamp 1626908933
transform 1 0 4368 0 1 19795
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2381
timestamp 1626908933
transform 1 0 4368 0 1 19795
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_128
timestamp 1626908933
transform -1 0 4512 0 -1 19980
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_59
timestamp 1626908933
transform -1 0 4512 0 -1 19980
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_279
timestamp 1626908933
transform 1 0 4512 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1270
timestamp 1626908933
transform 1 0 4512 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_444
timestamp 1626908933
transform 1 0 4752 0 1 19795
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2411
timestamp 1626908933
transform 1 0 4752 0 1 19795
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1830
timestamp 1626908933
transform 1 0 4560 0 1 19573
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3765
timestamp 1626908933
transform 1 0 4560 0 1 19573
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_273
timestamp 1626908933
transform 1 0 5300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_921
timestamp 1626908933
transform 1 0 5300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_273
timestamp 1626908933
transform 1 0 5300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_921
timestamp 1626908933
transform 1 0 5300 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_618
timestamp 1626908933
transform 1 0 4608 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1340
timestamp 1626908933
transform 1 0 4608 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_11
timestamp 1626908933
transform -1 0 5952 0 -1 19980
box -38 -49 614 715
use sky130_fd_sc_hs__o22ai_1  sky130_fd_sc_hs__o22ai_1_5
timestamp 1626908933
transform -1 0 5952 0 -1 19980
box -38 -49 614 715
use L1M1_PR  L1M1_PR_3176
timestamp 1626908933
transform 1 0 5424 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1241
timestamp 1626908933
transform 1 0 5424 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_399
timestamp 1626908933
transform 1 0 5808 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2366
timestamp 1626908933
transform 1 0 5808 0 1 19203
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1239
timestamp 1626908933
transform 1 0 5712 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3174
timestamp 1626908933
transform 1 0 5712 0 1 19425
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2477
timestamp 1626908933
transform 1 0 5616 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_510
timestamp 1626908933
transform 1 0 5616 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3819
timestamp 1626908933
transform 1 0 6192 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1852
timestamp 1626908933
transform 1 0 6192 0 1 19573
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2440
timestamp 1626908933
transform 1 0 5616 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_505
timestamp 1626908933
transform 1 0 5616 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2378
timestamp 1626908933
transform 1 0 5712 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_443
timestamp 1626908933
transform 1 0 5712 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3178
timestamp 1626908933
transform 1 0 5904 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1243
timestamp 1626908933
transform 1 0 5904 0 1 19721
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3149
timestamp 1626908933
transform 1 0 5904 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1182
timestamp 1626908933
transform 1 0 5904 0 1 19721
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_592
timestamp 1626908933
transform 1 0 5952 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1314
timestamp 1626908933
transform 1 0 5952 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_884
timestamp 1626908933
transform 1 0 6720 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1875
timestamp 1626908933
transform 1 0 6720 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1851
timestamp 1626908933
transform 1 0 6768 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3818
timestamp 1626908933
transform 1 0 6768 0 1 19573
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1828
timestamp 1626908933
transform 1 0 6768 0 1 19573
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3763
timestamp 1626908933
transform 1 0 6768 0 1 19573
box -29 -23 29 23
use M1M2_PR  M1M2_PR_443
timestamp 1626908933
transform 1 0 7152 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_450
timestamp 1626908933
transform 1 0 6960 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2410
timestamp 1626908933
transform 1 0 7152 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2417
timestamp 1626908933
transform 1 0 6960 0 1 19721
box -32 -32 32 32
use L1M1_PR  L1M1_PR_441
timestamp 1626908933
transform 1 0 7152 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_450
timestamp 1626908933
transform 1 0 7056 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2376
timestamp 1626908933
transform 1 0 7152 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2385
timestamp 1626908933
transform 1 0 7056 0 1 19721
box -29 -23 29 23
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_0
timestamp 1626908933
transform 1 0 6816 0 -1 19980
box -38 -49 710 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_5
timestamp 1626908933
transform 1 0 6816 0 -1 19980
box -38 -49 710 715
use L1M1_PR  L1M1_PR_2377
timestamp 1626908933
transform 1 0 7248 0 1 19795
box -29 -23 29 23
use L1M1_PR  L1M1_PR_442
timestamp 1626908933
transform 1 0 7248 0 1 19795
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_897
timestamp 1626908933
transform 1 0 7700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_249
timestamp 1626908933
transform 1 0 7700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_897
timestamp 1626908933
transform 1 0 7700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_249
timestamp 1626908933
transform 1 0 7700 0 1 19314
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2383
timestamp 1626908933
transform 1 0 7440 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_448
timestamp 1626908933
transform 1 0 7440 0 1 19721
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_502
timestamp 1626908933
transform 1 0 7488 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_145
timestamp 1626908933
transform 1 0 7488 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_746
timestamp 1626908933
transform 1 0 7584 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_145
timestamp 1626908933
transform 1 0 7584 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_278
timestamp 1626908933
transform 1 0 7776 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1269
timestamp 1626908933
transform 1 0 7776 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_554
timestamp 1626908933
transform 1 0 7872 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1276
timestamp 1626908933
transform 1 0 7872 0 -1 19980
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2414
timestamp 1626908933
transform 1 0 8112 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_447
timestamp 1626908933
transform 1 0 8112 0 1 19721
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_277
timestamp 1626908933
transform 1 0 8640 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1268
timestamp 1626908933
transform 1 0 8640 0 -1 19980
box -38 -49 134 715
use L1M1_PR  L1M1_PR_440
timestamp 1626908933
transform 1 0 8880 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_491
timestamp 1626908933
transform 1 0 8784 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2375
timestamp 1626908933
transform 1 0 8880 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2426
timestamp 1626908933
transform 1 0 8784 0 1 19721
box -29 -23 29 23
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_1
timestamp 1626908933
transform 1 0 8736 0 -1 19980
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_14
timestamp 1626908933
transform 1 0 8736 0 -1 19980
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2210
timestamp 1626908933
transform 1 0 9072 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2179
timestamp 1626908933
transform 1 0 8976 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_275
timestamp 1626908933
transform 1 0 9072 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_244
timestamp 1626908933
transform 1 0 8976 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2191
timestamp 1626908933
transform 1 0 8976 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_224
timestamp 1626908933
transform 1 0 8976 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2415
timestamp 1626908933
transform 1 0 9360 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_480
timestamp 1626908933
transform 1 0 9360 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2218
timestamp 1626908933
transform 1 0 9552 0 1 19499
box -32 -32 32 32
use M1M2_PR  M1M2_PR_251
timestamp 1626908933
transform 1 0 9552 0 1 19499
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1267
timestamp 1626908933
transform 1 0 9312 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_276
timestamp 1626908933
transform 1 0 9312 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1033
timestamp 1626908933
transform 1 0 9408 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_435
timestamp 1626908933
transform 1 0 9408 0 -1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_494
timestamp 1626908933
transform 1 0 9648 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2461
timestamp 1626908933
transform 1 0 9648 0 1 19869
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_225
timestamp 1626908933
transform 1 0 10100 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_873
timestamp 1626908933
transform 1 0 10100 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_225
timestamp 1626908933
transform 1 0 10100 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_873
timestamp 1626908933
transform 1 0 10100 0 1 19314
box -100 -49 100 49
use M1M2_PR  M1M2_PR_482
timestamp 1626908933
transform 1 0 9840 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2449
timestamp 1626908933
transform 1 0 9840 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1730
timestamp 1626908933
transform 1 0 10032 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3697
timestamp 1626908933
transform 1 0 10032 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_242
timestamp 1626908933
transform 1 0 9936 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2177
timestamp 1626908933
transform 1 0 9936 0 1 19721
box -29 -23 29 23
use M1M2_PR  M1M2_PR_490
timestamp 1626908933
transform 1 0 10512 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2457
timestamp 1626908933
transform 1 0 10512 0 1 19869
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_50
timestamp 1626908933
transform -1 0 12480 0 -1 19980
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_4
timestamp 1626908933
transform -1 0 12480 0 -1 19980
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_2365
timestamp 1626908933
transform 1 0 11856 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_398
timestamp 1626908933
transform 1 0 11856 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1021
timestamp 1626908933
transform 1 0 12048 0 1 19129
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2988
timestamp 1626908933
transform 1 0 12048 0 1 19129
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1711
timestamp 1626908933
transform 1 0 12048 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3646
timestamp 1626908933
transform 1 0 12048 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1622
timestamp 1626908933
transform 1 0 12336 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3589
timestamp 1626908933
transform 1 0 12336 0 1 19721
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1672
timestamp 1626908933
transform 1 0 12432 0 1 19573
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3607
timestamp 1626908933
transform 1 0 12432 0 1 19573
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_201
timestamp 1626908933
transform 1 0 12500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_849
timestamp 1626908933
transform 1 0 12500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_201
timestamp 1626908933
transform 1 0 12500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_849
timestamp 1626908933
transform 1 0 12500 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_144
timestamp 1626908933
transform 1 0 12480 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_501
timestamp 1626908933
transform 1 0 12480 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_144
timestamp 1626908933
transform 1 0 12576 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_745
timestamp 1626908933
transform 1 0 12576 0 -1 19980
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1671
timestamp 1626908933
transform 1 0 12528 0 1 19203
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3606
timestamp 1626908933
transform 1 0 12528 0 1 19203
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1582
timestamp 1626908933
transform 1 0 12720 0 1 19499
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1583
timestamp 1626908933
transform 1 0 12720 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1617
timestamp 1626908933
transform 1 0 12720 0 1 19795
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3549
timestamp 1626908933
transform 1 0 12720 0 1 19499
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3550
timestamp 1626908933
transform 1 0 12720 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3584
timestamp 1626908933
transform 1 0 12720 0 1 19795
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_109
timestamp 1626908933
transform 1 0 13536 0 -1 19980
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_47
timestamp 1626908933
transform 1 0 13536 0 -1 19980
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3057
timestamp 1626908933
transform 1 0 13488 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1122
timestamp 1626908933
transform 1 0 13488 0 1 19425
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3022
timestamp 1626908933
transform 1 0 13488 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1055
timestamp 1626908933
transform 1 0 13488 0 1 19425
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1181
timestamp 1626908933
transform 1 0 12768 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_459
timestamp 1626908933
transform 1 0 12768 0 -1 19980
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3062
timestamp 1626908933
transform 1 0 13776 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1127
timestamp 1626908933
transform 1 0 13776 0 1 19425
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1266
timestamp 1626908933
transform 1 0 13824 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_275
timestamp 1626908933
transform 1 0 13824 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1058
timestamp 1626908933
transform 1 0 14256 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3025
timestamp 1626908933
transform 1 0 14256 0 1 19425
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_177
timestamp 1626908933
transform 1 0 14900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_825
timestamp 1626908933
transform 1 0 14900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_177
timestamp 1626908933
transform 1 0 14900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_825
timestamp 1626908933
transform 1 0 14900 0 1 19314
box -100 -49 100 49
use M1M2_PR  M1M2_PR_249
timestamp 1626908933
transform 1 0 14640 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1053
timestamp 1626908933
transform 1 0 14064 0 1 19499
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2216
timestamp 1626908933
transform 1 0 14640 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3020
timestamp 1626908933
transform 1 0 14064 0 1 19499
box -32 -32 32 32
use L1M1_PR  L1M1_PR_272
timestamp 1626908933
transform 1 0 14736 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1120
timestamp 1626908933
transform 1 0 13872 0 1 19499
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2207
timestamp 1626908933
transform 1 0 14736 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3055
timestamp 1626908933
transform 1 0 13872 0 1 19499
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_428
timestamp 1626908933
transform 1 0 13920 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1150
timestamp 1626908933
transform 1 0 13920 0 -1 19980
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3591
timestamp 1626908933
transform 1 0 16368 0 1 19203
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1656
timestamp 1626908933
transform 1 0 16368 0 1 19203
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3677
timestamp 1626908933
transform 1 0 16464 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1710
timestamp 1626908933
transform 1 0 16464 0 1 19573
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_63
timestamp 1626908933
transform -1 0 17376 0 -1 19980
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_17
timestamp 1626908933
transform -1 0 17376 0 -1 19980
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_1701
timestamp 1626908933
transform 1 0 16944 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3636
timestamp 1626908933
transform 1 0 16944 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1566
timestamp 1626908933
transform 1 0 17040 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1567
timestamp 1626908933
transform 1 0 17040 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3533
timestamp 1626908933
transform 1 0 17040 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3534
timestamp 1626908933
transform 1 0 17040 0 1 19203
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_885
timestamp 1626908933
transform 1 0 17376 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1876
timestamp 1626908933
transform 1 0 17376 0 -1 19980
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1655
timestamp 1626908933
transform 1 0 17328 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3590
timestamp 1626908933
transform 1 0 17328 0 1 19647
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_153
timestamp 1626908933
transform 1 0 17300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_801
timestamp 1626908933
transform 1 0 17300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_153
timestamp 1626908933
transform 1 0 17300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_801
timestamp 1626908933
transform 1 0 17300 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_143
timestamp 1626908933
transform 1 0 17472 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_500
timestamp 1626908933
transform 1 0 17472 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_274
timestamp 1626908933
transform 1 0 17568 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1265
timestamp 1626908933
transform 1 0 17568 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_273
timestamp 1626908933
transform 1 0 18048 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1264
timestamp 1626908933
transform 1 0 18048 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_354
timestamp 1626908933
transform 1 0 18144 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1076
timestamp 1626908933
transform 1 0 18144 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_266
timestamp 1626908933
transform 1 0 17664 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_864
timestamp 1626908933
transform 1 0 17664 0 -1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3666
timestamp 1626908933
transform 1 0 18768 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1699
timestamp 1626908933
transform 1 0 18768 0 1 19573
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1263
timestamp 1626908933
transform 1 0 18912 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_272
timestamp 1626908933
transform 1 0 18912 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_837
timestamp 1626908933
transform 1 0 19008 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_239
timestamp 1626908933
transform 1 0 19008 0 -1 19980
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_777
timestamp 1626908933
transform 1 0 19700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_129
timestamp 1626908933
transform 1 0 19700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_777
timestamp 1626908933
transform 1 0 19700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_129
timestamp 1626908933
transform 1 0 19700 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1262
timestamp 1626908933
transform 1 0 20160 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_271
timestamp 1626908933
transform 1 0 20160 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1047
timestamp 1626908933
transform 1 0 19392 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_325
timestamp 1626908933
transform 1 0 19392 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_814
timestamp 1626908933
transform 1 0 20256 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_216
timestamp 1626908933
transform 1 0 20256 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1020
timestamp 1626908933
transform 1 0 20640 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_298
timestamp 1626908933
transform 1 0 20640 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1261
timestamp 1626908933
transform 1 0 21600 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_270
timestamp 1626908933
transform 1 0 21600 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_744
timestamp 1626908933
transform 1 0 21408 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_143
timestamp 1626908933
transform 1 0 21408 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_993
timestamp 1626908933
transform 1 0 21696 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_271
timestamp 1626908933
transform 1 0 21696 0 -1 19980
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_753
timestamp 1626908933
transform 1 0 22100 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_105
timestamp 1626908933
transform 1 0 22100 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_753
timestamp 1626908933
transform 1 0 22100 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_105
timestamp 1626908933
transform 1 0 22100 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_142
timestamp 1626908933
transform 1 0 22464 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_499
timestamp 1626908933
transform 1 0 22464 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_11
timestamp 1626908933
transform 1 0 22416 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1978
timestamp 1626908933
transform 1 0 22416 0 1 19203
box -32 -32 32 32
use L1M1_PR  L1M1_PR_13
timestamp 1626908933
transform 1 0 22320 0 1 19203
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1948
timestamp 1626908933
transform 1 0 22320 0 1 19203
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_525
timestamp 1626908933
transform 1 0 23328 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1126
timestamp 1626908933
transform 1 0 23328 0 -1 19980
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1341
timestamp 1626908933
transform 1 0 23088 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3308
timestamp 1626908933
transform 1 0 23088 0 1 19721
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_246
timestamp 1626908933
transform 1 0 22560 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_968
timestamp 1626908933
transform 1 0 22560 0 -1 19980
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3415
timestamp 1626908933
transform 1 0 23952 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1480
timestamp 1626908933
transform 1 0 23952 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3446
timestamp 1626908933
transform 1 0 23760 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3356
timestamp 1626908933
transform 1 0 23568 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1511
timestamp 1626908933
transform 1 0 23760 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1421
timestamp 1626908933
transform 1 0 23568 0 1 19721
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3394
timestamp 1626908933
transform 1 0 23664 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1427
timestamp 1626908933
transform 1 0 23664 0 1 19721
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_31
timestamp 1626908933
transform 1 0 23520 0 -1 19980
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_6
timestamp 1626908933
transform 1 0 23520 0 -1 19980
box -38 -49 518 715
use M1M2_PR  M1M2_PR_2335
timestamp 1626908933
transform 1 0 24336 0 1 19203
box -32 -32 32 32
use M1M2_PR  M1M2_PR_368
timestamp 1626908933
transform 1 0 24336 0 1 19203
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_729
timestamp 1626908933
transform 1 0 24500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_81
timestamp 1626908933
transform 1 0 24500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_729
timestamp 1626908933
transform 1 0 24500 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_81
timestamp 1626908933
transform 1 0 24500 0 1 19314
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3363
timestamp 1626908933
transform 1 0 24240 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1396
timestamp 1626908933
transform 1 0 24240 0 1 19425
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3425
timestamp 1626908933
transform 1 0 24816 0 1 19721
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1490
timestamp 1626908933
transform 1 0 24816 0 1 19721
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_202
timestamp 1626908933
transform 1 0 24000 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_924
timestamp 1626908933
transform 1 0 24000 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_55
timestamp 1626908933
transform 1 0 24768 0 -1 19980
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_9
timestamp 1626908933
transform 1 0 24768 0 -1 19980
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3395
timestamp 1626908933
transform 1 0 25200 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1460
timestamp 1626908933
transform 1 0 25200 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3346
timestamp 1626908933
transform 1 0 25488 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1379
timestamp 1626908933
transform 1 0 25488 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3374
timestamp 1626908933
transform 1 0 25872 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1407
timestamp 1626908933
transform 1 0 25872 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2349
timestamp 1626908933
transform 1 0 26544 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_382
timestamp 1626908933
transform 1 0 26544 0 1 19573
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_705
timestamp 1626908933
transform 1 0 26900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_57
timestamp 1626908933
transform 1 0 26900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_705
timestamp 1626908933
transform 1 0 26900 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_57
timestamp 1626908933
transform 1 0 26900 0 1 19314
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2326
timestamp 1626908933
transform 1 0 27312 0 1 19203
box -29 -23 29 23
use L1M1_PR  L1M1_PR_391
timestamp 1626908933
transform 1 0 27312 0 1 19203
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_743
timestamp 1626908933
transform 1 0 27552 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_142
timestamp 1626908933
transform 1 0 27552 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_498
timestamp 1626908933
transform 1 0 27456 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_141
timestamp 1626908933
transform 1 0 27456 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2321
timestamp 1626908933
transform 1 0 27696 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_354
timestamp 1626908933
transform 1 0 27696 0 1 19869
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_846
timestamp 1626908933
transform 1 0 27744 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_124
timestamp 1626908933
transform 1 0 27744 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_269
timestamp 1626908933
transform 1 0 28896 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1260
timestamp 1626908933
transform 1 0 28896 0 -1 19980
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_33
timestamp 1626908933
transform 1 0 29300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_681
timestamp 1626908933
transform 1 0 29300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_33
timestamp 1626908933
transform 1 0 29300 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_681
timestamp 1626908933
transform 1 0 29300 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_89
timestamp 1626908933
transform 1 0 28992 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_811
timestamp 1626908933
transform 1 0 28992 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_61
timestamp 1626908933
transform 1 0 28512 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_659
timestamp 1626908933
transform 1 0 28512 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_742
timestamp 1626908933
transform 1 0 29760 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_141
timestamp 1626908933
transform 1 0 29760 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_627
timestamp 1626908933
transform 1 0 29952 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_29
timestamp 1626908933
transform 1 0 29952 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_21
timestamp 1626908933
transform 1 0 30336 0 -1 19980
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_6
timestamp 1626908933
transform 1 0 30336 0 -1 19980
box -38 -49 710 715
use L1M1_PR  L1M1_PR_1815
timestamp 1626908933
transform 1 0 30480 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3750
timestamp 1626908933
transform 1 0 30480 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_411
timestamp 1626908933
transform 1 0 30672 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1882
timestamp 1626908933
transform 1 0 30768 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2378
timestamp 1626908933
transform 1 0 30672 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3849
timestamp 1626908933
transform 1 0 30768 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_404
timestamp 1626908933
transform 1 0 30672 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1857
timestamp 1626908933
transform 1 0 30768 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2339
timestamp 1626908933
transform 1 0 30672 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3792
timestamp 1626908933
transform 1 0 30768 0 1 19647
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_268
timestamp 1626908933
transform 1 0 31008 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1259
timestamp 1626908933
transform 1 0 31008 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_403
timestamp 1626908933
transform 1 0 30960 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1825
timestamp 1626908933
transform 1 0 31056 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2370
timestamp 1626908933
transform 1 0 30960 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3792
timestamp 1626908933
transform 1 0 31056 0 1 19721
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1796
timestamp 1626908933
transform 1 0 30960 0 1 19425
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3731
timestamp 1626908933
transform 1 0 30960 0 1 19425
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_6
timestamp 1626908933
transform 1 0 31104 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_604
timestamp 1626908933
transform 1 0 31104 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_267
timestamp 1626908933
transform 1 0 31488 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1258
timestamp 1626908933
transform 1 0 31488 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1789
timestamp 1626908933
transform 1 0 31344 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3756
timestamp 1626908933
transform 1 0 31344 0 1 19425
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_140
timestamp 1626908933
transform 1 0 31680 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_497
timestamp 1626908933
transform 1 0 31680 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_886
timestamp 1626908933
transform 1 0 31584 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1877
timestamp 1626908933
transform 1 0 31584 0 -1 19980
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_9
timestamp 1626908933
transform 1 0 31700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_657
timestamp 1626908933
transform 1 0 31700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_9
timestamp 1626908933
transform 1 0 31700 0 1 19314
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_657
timestamp 1626908933
transform 1 0 31700 0 1 19314
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_526
timestamp 1626908933
transform 1 0 31776 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1127
timestamp 1626908933
transform 1 0 31776 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1878
timestamp 1626908933
transform 1 0 31968 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_887
timestamp 1626908933
transform 1 0 31968 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3830
timestamp 1626908933
transform 1 0 48 0 1 20165
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1863
timestamp 1626908933
transform 1 0 48 0 1 20165
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1879
timestamp 1626908933
transform 1 0 192 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_888
timestamp 1626908933
transform 1 0 192 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3840
timestamp 1626908933
transform 1 0 240 0 1 20461
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1873
timestamp 1626908933
transform 1 0 240 0 1 20461
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_496
timestamp 1626908933
transform 1 0 288 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_139
timestamp 1626908933
transform 1 0 288 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1128
timestamp 1626908933
transform 1 0 0 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_736
timestamp 1626908933
transform 1 0 0 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_527
timestamp 1626908933
transform 1 0 0 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_135
timestamp 1626908933
transform 1 0 0 0 -1 21312
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_320
timestamp 1626908933
transform 1 0 500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_968
timestamp 1626908933
transform 1 0 500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_320
timestamp 1626908933
transform 1 0 500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_968
timestamp 1626908933
transform 1 0 500 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_694
timestamp 1626908933
transform 1 0 384 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_708
timestamp 1626908933
transform 1 0 192 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1416
timestamp 1626908933
transform 1 0 384 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1430
timestamp 1626908933
transform 1 0 192 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_256
timestamp 1626908933
transform 1 0 960 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1247
timestamp 1626908933
transform 1 0 960 0 -1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1541
timestamp 1626908933
transform 1 0 1200 0 1 20535
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3508
timestamp 1626908933
transform 1 0 1200 0 1 20535
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1627
timestamp 1626908933
transform 1 0 1200 0 1 20535
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3562
timestamp 1626908933
transform 1 0 1200 0 1 20535
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1281
timestamp 1626908933
transform 1 0 1700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_633
timestamp 1626908933
transform 1 0 1700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1281
timestamp 1626908933
transform 1 0 1700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_633
timestamp 1626908933
transform 1 0 1700 0 1 19980
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2978
timestamp 1626908933
transform 1 0 1392 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1043
timestamp 1626908933
transform 1 0 1392 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2948
timestamp 1626908933
transform 1 0 1392 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_981
timestamp 1626908933
transform 1 0 1392 0 1 20313
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2262
timestamp 1626908933
transform 1 0 1680 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_327
timestamp 1626908933
transform 1 0 1680 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3138
timestamp 1626908933
transform 1 0 1584 0 1 20535
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1203
timestamp 1626908933
transform 1 0 1584 0 1 20535
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3100
timestamp 1626908933
transform 1 0 1584 0 1 20535
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1133
timestamp 1626908933
transform 1 0 1584 0 1 20535
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_674
timestamp 1626908933
transform 1 0 1440 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1396
timestamp 1626908933
transform 1 0 1440 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_570
timestamp 1626908933
transform 1 0 1056 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1168
timestamp 1626908933
transform 1 0 1056 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_38
timestamp 1626908933
transform 1 0 1152 0 1 19980
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_77
timestamp 1626908933
transform 1 0 1152 0 1 19980
box -38 -49 614 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_132
timestamp 1626908933
transform 1 0 2496 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_489
timestamp 1626908933
transform 1 0 2496 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_530
timestamp 1626908933
transform 1 0 2304 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1131
timestamp 1626908933
transform 1 0 2304 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_255
timestamp 1626908933
transform 1 0 2208 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1246
timestamp 1626908933
transform 1 0 2208 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_661
timestamp 1626908933
transform 1 0 2112 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1383
timestamp 1626908933
transform 1 0 2112 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_554
timestamp 1626908933
transform 1 0 1728 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1152
timestamp 1626908933
transform 1 0 1728 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1144
timestamp 1626908933
transform 1 0 2592 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_546
timestamp 1626908933
transform 1 0 2592 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_36
timestamp 1626908933
transform 1 0 2976 0 -1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_97
timestamp 1626908933
transform 1 0 2976 0 -1 21312
box -38 -49 326 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_296
timestamp 1626908933
transform 1 0 2900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_944
timestamp 1626908933
transform 1 0 2900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_296
timestamp 1626908933
transform 1 0 2900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_944
timestamp 1626908933
transform 1 0 2900 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_254
timestamp 1626908933
transform 1 0 3264 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1245
timestamp 1626908933
transform 1 0 3264 0 -1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_303
timestamp 1626908933
transform 1 0 3312 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2270
timestamp 1626908933
transform 1 0 3312 0 1 20313
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_642
timestamp 1626908933
transform 1 0 3360 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_643
timestamp 1626908933
transform 1 0 3264 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1364
timestamp 1626908933
transform 1 0 3360 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1365
timestamp 1626908933
transform 1 0 3264 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_543
timestamp 1626908933
transform 1 0 2880 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1141
timestamp 1626908933
transform 1 0 2880 0 1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1860
timestamp 1626908933
transform 1 0 3984 0 1 20165
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3827
timestamp 1626908933
transform 1 0 3984 0 1 20165
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1837
timestamp 1626908933
transform 1 0 3984 0 1 20165
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3772
timestamp 1626908933
transform 1 0 3984 0 1 20165
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1257
timestamp 1626908933
transform 1 0 4100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_609
timestamp 1626908933
transform 1 0 4100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1257
timestamp 1626908933
transform 1 0 4100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_609
timestamp 1626908933
transform 1 0 4100 0 1 19980
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3782
timestamp 1626908933
transform 1 0 4176 0 1 20461
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1847
timestamp 1626908933
transform 1 0 4176 0 1 20461
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3839
timestamp 1626908933
transform 1 0 4176 0 1 20461
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1872
timestamp 1626908933
transform 1 0 4176 0 1 20461
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_735
timestamp 1626908933
transform 1 0 4416 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_134
timestamp 1626908933
transform 1 0 4416 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_112
timestamp 1626908933
transform -1 0 4416 0 -1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_51
timestamp 1626908933
transform -1 0 4416 0 -1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_3
timestamp 1626908933
transform 1 0 4032 0 1 19980
box -38 -49 614 715
use sky130_fd_sc_hs__o31ai_1  sky130_fd_sc_hs__o31ai_1_7
timestamp 1626908933
transform 1 0 4032 0 1 19980
box -38 -49 614 715
use M1M2_PR  M1M2_PR_504
timestamp 1626908933
transform 1 0 4752 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2471
timestamp 1626908933
transform 1 0 4752 0 1 20313
box -32 -32 32 32
use L1M1_PR  L1M1_PR_498
timestamp 1626908933
transform 1 0 4656 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1238
timestamp 1626908933
transform 1 0 4560 0 1 20091
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1271
timestamp 1626908933
transform 1 0 4464 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2433
timestamp 1626908933
transform 1 0 4656 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3173
timestamp 1626908933
transform 1 0 4560 0 1 20091
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3206
timestamp 1626908933
transform 1 0 4464 0 1 20313
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_138
timestamp 1626908933
transform 1 0 4992 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_495
timestamp 1626908933
transform 1 0 4992 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1176
timestamp 1626908933
transform 1 0 4944 0 1 20091
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3143
timestamp 1626908933
transform 1 0 4944 0 1 20091
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_272
timestamp 1626908933
transform 1 0 5300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_920
timestamp 1626908933
transform 1 0 5300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_272
timestamp 1626908933
transform 1 0 5300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_920
timestamp 1626908933
transform 1 0 5300 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_617
timestamp 1626908933
transform 1 0 4608 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1339
timestamp 1626908933
transform 1 0 4608 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_40
timestamp 1626908933
transform 1 0 4608 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_41
timestamp 1626908933
transform 1 0 5088 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_92
timestamp 1626908933
transform 1 0 4608 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_93
timestamp 1626908933
transform 1 0 5088 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2432
timestamp 1626908933
transform 1 0 5520 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_497
timestamp 1626908933
transform 1 0 5520 0 1 20313
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1884
timestamp 1626908933
transform 1 0 5376 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_893
timestamp 1626908933
transform 1 0 5376 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1129
timestamp 1626908933
transform 1 0 5472 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_528
timestamp 1626908933
transform 1 0 5472 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_113
timestamp 1626908933
transform 1 0 5472 0 -1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_52
timestamp 1626908933
transform 1 0 5472 0 -1 21312
box -38 -49 326 715
use M1M2_PR  M1M2_PR_2476
timestamp 1626908933
transform 1 0 5616 0 1 20165
box -32 -32 32 32
use M1M2_PR  M1M2_PR_509
timestamp 1626908933
transform 1 0 5616 0 1 20165
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1244
timestamp 1626908933
transform 1 0 5760 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_253
timestamp 1626908933
transform 1 0 5760 0 -1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2438
timestamp 1626908933
transform 1 0 5904 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2429
timestamp 1626908933
transform 1 0 6000 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_503
timestamp 1626908933
transform 1 0 5904 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_494
timestamp 1626908933
transform 1 0 6000 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2467
timestamp 1626908933
transform 1 0 6000 0 1 20091
box -32 -32 32 32
use M1M2_PR  M1M2_PR_500
timestamp 1626908933
transform 1 0 6000 0 1 20091
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2431
timestamp 1626908933
transform 1 0 6096 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2370
timestamp 1626908933
transform 1 0 6096 0 1 20387
box -29 -23 29 23
use L1M1_PR  L1M1_PR_496
timestamp 1626908933
transform 1 0 6096 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_435
timestamp 1626908933
transform 1 0 6096 0 1 20387
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_585
timestamp 1626908933
transform 1 0 6500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1233
timestamp 1626908933
transform 1 0 6500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_585
timestamp 1626908933
transform 1 0 6500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1233
timestamp 1626908933
transform 1 0 6500 0 1 19980
box -100 -49 100 49
use M1M2_PR  M1M2_PR_507
timestamp 1626908933
transform 1 0 6288 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2474
timestamp 1626908933
transform 1 0 6288 0 1 20239
box -32 -32 32 32
use L1M1_PR  L1M1_PR_501
timestamp 1626908933
transform 1 0 6288 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2436
timestamp 1626908933
transform 1 0 6288 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_247
timestamp 1626908933
transform 1 0 6672 0 1 20165
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2182
timestamp 1626908933
transform 1 0 6672 0 1 20165
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2406
timestamp 1626908933
transform 1 0 6576 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_439
timestamp 1626908933
transform 1 0 6576 0 1 20387
box -32 -32 32 32
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_13
timestamp 1626908933
transform -1 0 7200 0 -1 21312
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_0
timestamp 1626908933
transform -1 0 7200 0 -1 21312
box -38 -49 614 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_591
timestamp 1626908933
transform 1 0 5856 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1313
timestamp 1626908933
transform 1 0 5856 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_1
timestamp 1626908933
transform 1 0 5664 0 1 19980
box -38 -49 710 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_6
timestamp 1626908933
transform 1 0 5664 0 1 19980
box -38 -49 710 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_531
timestamp 1626908933
transform 1 0 7200 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1132
timestamp 1626908933
transform 1 0 7200 0 -1 21312
box -38 -49 230 715
use L1M1_PR  L1M1_PR_439
timestamp 1626908933
transform 1 0 7152 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2374
timestamp 1626908933
transform 1 0 7152 0 1 19869
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3600
timestamp 1626908933
transform 1 0 7536 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1633
timestamp 1626908933
transform 1 0 7536 0 1 20313
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1885
timestamp 1626908933
transform 1 0 7392 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_894
timestamp 1626908933
transform 1 0 7392 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_488
timestamp 1626908933
transform 1 0 7488 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_131
timestamp 1626908933
transform 1 0 7488 0 -1 21312
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_896
timestamp 1626908933
transform 1 0 7700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_248
timestamp 1626908933
transform 1 0 7700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_896
timestamp 1626908933
transform 1 0 7700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_248
timestamp 1626908933
transform 1 0 7700 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1063
timestamp 1626908933
transform 1 0 7584 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_465
timestamp 1626908933
transform 1 0 7584 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_532
timestamp 1626908933
transform 1 0 7968 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1133
timestamp 1626908933
transform 1 0 7968 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_895
timestamp 1626908933
transform 1 0 8160 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1886
timestamp 1626908933
transform 1 0 8160 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_60
timestamp 1626908933
transform 1 0 8256 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_122
timestamp 1626908933
transform 1 0 8256 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_73
timestamp 1626908933
transform -1 0 9024 0 1 19980
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_27
timestamp 1626908933
transform -1 0 9024 0 1 19980
box -38 -49 2726 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1209
timestamp 1626908933
transform 1 0 8900 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_561
timestamp 1626908933
transform 1 0 8900 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1209
timestamp 1626908933
transform 1 0 8900 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_561
timestamp 1626908933
transform 1 0 8900 0 1 19980
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2250
timestamp 1626908933
transform 1 0 8688 0 1 20165
box -32 -32 32 32
use M1M2_PR  M1M2_PR_283
timestamp 1626908933
transform 1 0 8688 0 1 20165
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2430
timestamp 1626908933
transform 1 0 9072 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_463
timestamp 1626908933
transform 1 0 9072 0 1 20239
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2399
timestamp 1626908933
transform 1 0 9264 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_464
timestamp 1626908933
transform 1 0 9264 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3170
timestamp 1626908933
transform 1 0 8304 0 1 20535
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1203
timestamp 1626908933
transform 1 0 8304 0 1 20535
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3648
timestamp 1626908933
transform 1 0 8592 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1713
timestamp 1626908933
transform 1 0 8592 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3605
timestamp 1626908933
transform 1 0 8976 0 1 20387
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1670
timestamp 1626908933
transform 1 0 8976 0 1 20387
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2398
timestamp 1626908933
transform 1 0 9072 0 1 20535
box -29 -23 29 23
use L1M1_PR  L1M1_PR_463
timestamp 1626908933
transform 1 0 9072 0 1 20535
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2429
timestamp 1626908933
transform 1 0 9072 0 1 20535
box -32 -32 32 32
use M1M2_PR  M1M2_PR_462
timestamp 1626908933
transform 1 0 9072 0 1 20535
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_16
timestamp 1626908933
transform 1 0 8640 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_39
timestamp 1626908933
transform 1 0 8640 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__a222o_1  sky130_fd_sc_hs__a222o_1_0
timestamp 1626908933
transform -1 0 9984 0 1 19980
box -38 -49 998 715
use sky130_fd_sc_hs__a222o_1  sky130_fd_sc_hs__a222o_1_1
timestamp 1626908933
transform -1 0 9984 0 1 19980
box -38 -49 998 715
use L1M1_PR  L1M1_PR_2424
timestamp 1626908933
transform 1 0 9648 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2240
timestamp 1626908933
transform 1 0 9360 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_489
timestamp 1626908933
transform 1 0 9648 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_305
timestamp 1626908933
transform 1 0 9360 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2460
timestamp 1626908933
transform 1 0 9648 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_493
timestamp 1626908933
transform 1 0 9648 0 1 20239
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2414
timestamp 1626908933
transform 1 0 9744 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2181
timestamp 1626908933
transform 1 0 9456 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_479
timestamp 1626908933
transform 1 0 9744 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_246
timestamp 1626908933
transform 1 0 9456 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2448
timestamp 1626908933
transform 1 0 9840 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2193
timestamp 1626908933
transform 1 0 9552 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_481
timestamp 1626908933
transform 1 0 9840 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_226
timestamp 1626908933
transform 1 0 9552 0 1 20313
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_62
timestamp 1626908933
transform -1 0 9792 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_0
timestamp 1626908933
transform -1 0 9792 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1030
timestamp 1626908933
transform 1 0 9792 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_432
timestamp 1626908933
transform 1 0 9792 0 -1 21312
box -38 -49 422 715
use L1M1_PR  L1M1_PR_278
timestamp 1626908933
transform 1 0 9936 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2213
timestamp 1626908933
transform 1 0 9936 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1729
timestamp 1626908933
transform 1 0 10032 0 1 20461
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3696
timestamp 1626908933
transform 1 0 10032 0 1 20461
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_224
timestamp 1626908933
transform 1 0 10100 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_872
timestamp 1626908933
transform 1 0 10100 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_224
timestamp 1626908933
transform 1 0 10100 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_872
timestamp 1626908933
transform 1 0 10100 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_137
timestamp 1626908933
transform 1 0 9984 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_494
timestamp 1626908933
transform 1 0 9984 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1134
timestamp 1626908933
transform 1 0 10176 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_533
timestamp 1626908933
transform 1 0 10176 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1018
timestamp 1626908933
transform 1 0 10080 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_420
timestamp 1626908933
transform 1 0 10080 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_113
timestamp 1626908933
transform 1 0 10368 0 -1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_44
timestamp 1626908933
transform 1 0 10368 0 -1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1243
timestamp 1626908933
transform 1 0 10848 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_252
timestamp 1626908933
transform 1 0 10848 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1233
timestamp 1626908933
transform 1 0 10464 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1216
timestamp 1626908933
transform 1 0 10944 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_511
timestamp 1626908933
transform 1 0 10464 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_494
timestamp 1626908933
transform 1 0 10944 0 -1 21312
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1185
timestamp 1626908933
transform 1 0 11300 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_537
timestamp 1626908933
transform 1 0 11300 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1185
timestamp 1626908933
transform 1 0 11300 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_537
timestamp 1626908933
transform 1 0 11300 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_741
timestamp 1626908933
transform 1 0 11232 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_140
timestamp 1626908933
transform 1 0 11232 0 1 19980
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3548
timestamp 1626908933
transform 1 0 11472 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1581
timestamp 1626908933
transform 1 0 11472 0 1 20387
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1257
timestamp 1626908933
transform 1 0 11424 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_266
timestamp 1626908933
transform 1 0 11424 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_103
timestamp 1626908933
transform -1 0 12096 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_41
timestamp 1626908933
transform -1 0 12096 0 -1 21312
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1565
timestamp 1626908933
transform 1 0 12144 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3532
timestamp 1626908933
transform 1 0 12144 0 1 20387
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1654
timestamp 1626908933
transform 1 0 12336 0 1 20387
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3589
timestamp 1626908933
transform 1 0 12336 0 1 20387
box -29 -23 29 23
use M1M2_PR  M1M2_PR_397
timestamp 1626908933
transform 1 0 11856 0 1 20461
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2364
timestamp 1626908933
transform 1 0 11856 0 1 20461
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_200
timestamp 1626908933
transform 1 0 12500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_848
timestamp 1626908933
transform 1 0 12500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_200
timestamp 1626908933
transform 1 0 12500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_848
timestamp 1626908933
transform 1 0 12500 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_976
timestamp 1626908933
transform 1 0 12096 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_378
timestamp 1626908933
transform 1 0 12096 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_480
timestamp 1626908933
transform 1 0 11520 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1202
timestamp 1626908933
transform 1 0 11520 0 1 19980
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3642
timestamp 1626908933
transform 1 0 12720 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1707
timestamp 1626908933
transform 1 0 12720 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3583
timestamp 1626908933
transform 1 0 12720 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1616
timestamp 1626908933
transform 1 0 12720 0 1 20313
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_487
timestamp 1626908933
transform 1 0 12480 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_130
timestamp 1626908933
transform 1 0 12480 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_107
timestamp 1626908933
transform -1 0 13344 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_45
timestamp 1626908933
transform -1 0 13344 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_958
timestamp 1626908933
transform 1 0 12576 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_360
timestamp 1626908933
transform 1 0 12576 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_734
timestamp 1626908933
transform 1 0 13344 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_133
timestamp 1626908933
transform 1 0 13344 0 -1 21312
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1161
timestamp 1626908933
transform 1 0 13700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_513
timestamp 1626908933
transform 1 0 13700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1161
timestamp 1626908933
transform 1 0 13700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_513
timestamp 1626908933
transform 1 0 13700 0 1 19980
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3690
timestamp 1626908933
transform 1 0 13488 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1723
timestamp 1626908933
transform 1 0 13488 0 1 20387
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1242
timestamp 1626908933
transform 1 0 13536 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_251
timestamp 1626908933
transform 1 0 13536 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_440
timestamp 1626908933
transform 1 0 13632 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1162
timestamp 1626908933
transform 1 0 13632 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_83
timestamp 1626908933
transform 1 0 12288 0 1 19980
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_37
timestamp 1626908933
transform 1 0 12288 0 1 19980
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1052
timestamp 1626908933
transform 1 0 14160 0 1 20091
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3019
timestamp 1626908933
transform 1 0 14160 0 1 20091
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_250
timestamp 1626908933
transform 1 0 14400 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_896
timestamp 1626908933
transform 1 0 14496 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1241
timestamp 1626908933
transform 1 0 14400 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1887
timestamp 1626908933
transform 1 0 14496 0 -1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_254
timestamp 1626908933
transform 1 0 14640 0 1 20165
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2221
timestamp 1626908933
transform 1 0 14640 0 1 20165
box -32 -32 32 32
use L1M1_PR  L1M1_PR_277
timestamp 1626908933
transform 1 0 14640 0 1 20165
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2212
timestamp 1626908933
transform 1 0 14640 0 1 20165
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_117
timestamp 1626908933
transform 1 0 14592 0 -1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_48
timestamp 1626908933
transform 1 0 14592 0 -1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_136
timestamp 1626908933
transform 1 0 14976 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_493
timestamp 1626908933
transform 1 0 14976 0 1 19980
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_176
timestamp 1626908933
transform 1 0 14900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_824
timestamp 1626908933
transform 1 0 14900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_176
timestamp 1626908933
transform 1 0 14900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_824
timestamp 1626908933
transform 1 0 14900 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_249
timestamp 1626908933
transform 1 0 15456 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_265
timestamp 1626908933
transform 1 0 15456 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1240
timestamp 1626908933
transform 1 0 15456 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1256
timestamp 1626908933
transform 1 0 15456 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_245
timestamp 1626908933
transform 1 0 15216 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2212
timestamp 1626908933
transform 1 0 15216 0 1 20239
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_317
timestamp 1626908933
transform 1 0 15072 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_318
timestamp 1626908933
transform 1 0 15072 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_915
timestamp 1626908933
transform 1 0 15072 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_916
timestamp 1626908933
transform 1 0 15072 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_264
timestamp 1626908933
transform 1 0 16320 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1255
timestamp 1626908933
transform 1 0 16320 0 1 19980
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_489
timestamp 1626908933
transform 1 0 16100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1137
timestamp 1626908933
transform 1 0 16100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_489
timestamp 1626908933
transform 1 0 16100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1137
timestamp 1626908933
transform 1 0 16100 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_406
timestamp 1626908933
transform 1 0 15552 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_407
timestamp 1626908933
transform 1 0 15552 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1128
timestamp 1626908933
transform 1 0 15552 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1129
timestamp 1626908933
transform 1 0 15552 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_295
timestamp 1626908933
transform 1 0 16320 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_893
timestamp 1626908933
transform 1 0 16320 0 -1 21312
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3053
timestamp 1626908933
transform 1 0 16560 0 1 20091
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2199
timestamp 1626908933
transform 1 0 16560 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1118
timestamp 1626908933
transform 1 0 16560 0 1 20091
box -29 -23 29 23
use L1M1_PR  L1M1_PR_264
timestamp 1626908933
transform 1 0 16560 0 1 20239
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1880
timestamp 1626908933
transform 1 0 16416 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_889
timestamp 1626908933
transform 1 0 16416 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_105
timestamp 1626908933
transform -1 0 16800 0 1 19980
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_44
timestamp 1626908933
transform -1 0 16800 0 1 19980
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3049
timestamp 1626908933
transform 1 0 16752 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1114
timestamp 1626908933
transform 1 0 16752 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3018
timestamp 1626908933
transform 1 0 16656 0 1 20091
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3016
timestamp 1626908933
transform 1 0 16848 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1051
timestamp 1626908933
transform 1 0 16656 0 1 20091
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1049
timestamp 1626908933
transform 1 0 16848 0 1 20239
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1254
timestamp 1626908933
transform 1 0 16800 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_263
timestamp 1626908933
transform 1 0 16800 0 1 19980
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_800
timestamp 1626908933
transform 1 0 17300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_152
timestamp 1626908933
transform 1 0 17300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_800
timestamp 1626908933
transform 1 0 17300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_152
timestamp 1626908933
transform 1 0 17300 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_885
timestamp 1626908933
transform 1 0 16896 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_287
timestamp 1626908933
transform 1 0 16896 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1950
timestamp 1626908933
transform 1 0 17424 0 1 20535
box -29 -23 29 23
use L1M1_PR  L1M1_PR_15
timestamp 1626908933
transform 1 0 17424 0 1 20535
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1980
timestamp 1626908933
transform 1 0 17520 0 1 20535
box -32 -32 32 32
use M1M2_PR  M1M2_PR_13
timestamp 1626908933
transform 1 0 17520 0 1 20535
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_486
timestamp 1626908933
transform 1 0 17472 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_129
timestamp 1626908933
transform 1 0 17472 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1888
timestamp 1626908933
transform 1 0 17760 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_897
timestamp 1626908933
transform 1 0 17760 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1135
timestamp 1626908933
transform 1 0 17568 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_534
timestamp 1626908933
transform 1 0 17568 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_378
timestamp 1626908933
transform 1 0 16704 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1100
timestamp 1626908933
transform 1 0 16704 0 -1 21312
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_465
timestamp 1626908933
transform 1 0 18500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1113
timestamp 1626908933
transform 1 0 18500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_465
timestamp 1626908933
transform 1 0 18500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1113
timestamp 1626908933
transform 1 0 18500 0 1 19980
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1537
timestamp 1626908933
transform 1 0 18192 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3504
timestamp 1626908933
transform 1 0 18192 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_396
timestamp 1626908933
transform 1 0 19056 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2363
timestamp 1626908933
transform 1 0 19056 0 1 20387
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1622
timestamp 1626908933
transform 1 0 19344 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3557
timestamp 1626908933
transform 1 0 19344 0 1 20239
box -29 -23 29 23
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_7
timestamp 1626908933
transform -1 0 19680 0 1 19980
box -38 -49 2438 715
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_4
timestamp 1626908933
transform 1 0 17856 0 -1 21312
box -38 -49 2438 715
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_3
timestamp 1626908933
transform -1 0 19680 0 1 19980
box -38 -49 2438 715
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_0
timestamp 1626908933
transform 1 0 17856 0 -1 21312
box -38 -49 2438 715
use L1M1_PR  L1M1_PR_2355
timestamp 1626908933
transform 1 0 19536 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_420
timestamp 1626908933
transform 1 0 19536 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2391
timestamp 1626908933
transform 1 0 19536 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_424
timestamp 1626908933
transform 1 0 19536 0 1 20239
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_776
timestamp 1626908933
transform 1 0 19700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_128
timestamp 1626908933
transform 1 0 19700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_776
timestamp 1626908933
transform 1 0 19700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_128
timestamp 1626908933
transform 1 0 19700 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1881
timestamp 1626908933
transform 1 0 19872 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_890
timestamp 1626908933
transform 1 0 19872 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1130
timestamp 1626908933
transform 1 0 19680 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_529
timestamp 1626908933
transform 1 0 19680 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_492
timestamp 1626908933
transform 1 0 19968 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_135
timestamp 1626908933
transform 1 0 19968 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3281
timestamp 1626908933
transform 1 0 20112 0 1 20535
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1314
timestamp 1626908933
transform 1 0 20112 0 1 20535
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_733
timestamp 1626908933
transform 1 0 20256 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_132
timestamp 1626908933
transform 1 0 20256 0 -1 21312
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3500
timestamp 1626908933
transform 1 0 20400 0 1 20091
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1533
timestamp 1626908933
transform 1 0 20400 0 1 20091
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1239
timestamp 1626908933
transform 1 0 20448 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_248
timestamp 1626908933
transform 1 0 20448 0 -1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3328
timestamp 1626908933
transform 1 0 20592 0 1 20535
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1393
timestamp 1626908933
transform 1 0 20592 0 1 20535
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_297
timestamp 1626908933
transform 1 0 20544 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1019
timestamp 1626908933
transform 1 0 20544 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_0
timestamp 1626908933
transform 1 0 21312 0 -1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_61
timestamp 1626908933
transform 1 0 21312 0 -1 21312
box -38 -49 326 715
use M1M2_PR  M1M2_PR_391
timestamp 1626908933
transform 1 0 21264 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2358
timestamp 1626908933
transform 1 0 21264 0 1 20313
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_441
timestamp 1626908933
transform 1 0 20900 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1089
timestamp 1626908933
transform 1 0 20900 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_441
timestamp 1626908933
transform 1 0 20900 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1089
timestamp 1626908933
transform 1 0 20900 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_247
timestamp 1626908933
transform 1 0 21600 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1238
timestamp 1626908933
transform 1 0 21600 0 -1 21312
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_104
timestamp 1626908933
transform 1 0 22100 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_752
timestamp 1626908933
transform 1 0 22100 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_104
timestamp 1626908933
transform 1 0 22100 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_752
timestamp 1626908933
transform 1 0 22100 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_270
timestamp 1626908933
transform 1 0 21696 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_992
timestamp 1626908933
transform 1 0 21696 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__dfsbp_2  sky130_fd_sc_hs__dfsbp_2_1
timestamp 1626908933
transform -1 0 22656 0 1 19980
box -38 -49 2630 715
use sky130_fd_sc_hs__dfsbp_2  sky130_fd_sc_hs__dfsbp_2_0
timestamp 1626908933
transform -1 0 22656 0 1 19980
box -38 -49 2630 715
use L1M1_PR  L1M1_PR_3554
timestamp 1626908933
transform 1 0 22320 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1619
timestamp 1626908933
transform 1 0 22320 0 1 20239
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1977
timestamp 1626908933
transform 1 0 22416 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_10
timestamp 1626908933
transform 1 0 22416 0 1 20239
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_485
timestamp 1626908933
transform 1 0 22464 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_128
timestamp 1626908933
transform 1 0 22464 0 -1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1947
timestamp 1626908933
transform 1 0 22512 0 1 20239
box -29 -23 29 23
use L1M1_PR  L1M1_PR_12
timestamp 1626908933
transform 1 0 22512 0 1 20239
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_740
timestamp 1626908933
transform 1 0 22656 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_139
timestamp 1626908933
transform 1 0 22656 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_769
timestamp 1626908933
transform 1 0 22560 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_171
timestamp 1626908933
transform 1 0 22560 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_172
timestamp 1626908933
transform 1 0 22848 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_770
timestamp 1626908933
transform 1 0 22848 0 1 19980
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_417
timestamp 1626908933
transform 1 0 23300 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1065
timestamp 1626908933
transform 1 0 23300 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_417
timestamp 1626908933
transform 1 0 23300 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1065
timestamp 1626908933
transform 1 0 23300 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_232
timestamp 1626908933
transform 1 0 23232 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_954
timestamp 1626908933
transform 1 0 23232 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_138
timestamp 1626908933
transform 1 0 24000 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_739
timestamp 1626908933
transform 1 0 24000 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_132
timestamp 1626908933
transform 1 0 24768 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_730
timestamp 1626908933
transform 1 0 24768 0 -1 21312
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_80
timestamp 1626908933
transform 1 0 24500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_728
timestamp 1626908933
transform 1 0 24500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_80
timestamp 1626908933
transform 1 0 24500 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_728
timestamp 1626908933
transform 1 0 24500 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_201
timestamp 1626908933
transform 1 0 24192 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_923
timestamp 1626908933
transform 1 0 24192 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_12
timestamp 1626908933
transform -1 0 24768 0 -1 21312
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_0
timestamp 1626908933
transform -1 0 24768 0 -1 21312
box -38 -49 1862 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_134
timestamp 1626908933
transform 1 0 24960 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_491
timestamp 1626908933
transform 1 0 24960 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_262
timestamp 1626908933
transform 1 0 25056 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1253
timestamp 1626908933
transform 1 0 25056 0 1 19980
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1041
timestamp 1626908933
transform 1 0 25700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_393
timestamp 1626908933
transform 1 0 25700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1041
timestamp 1626908933
transform 1 0 25700 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_393
timestamp 1626908933
transform 1 0 25700 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_738
timestamp 1626908933
transform 1 0 25920 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_137
timestamp 1626908933
transform 1 0 25920 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_39
timestamp 1626908933
transform -1 0 26400 0 -1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_14
timestamp 1626908933
transform -1 0 26400 0 -1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_702
timestamp 1626908933
transform 1 0 26112 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_104
timestamp 1626908933
transform 1 0 26112 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_182
timestamp 1626908933
transform 1 0 25152 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_183
timestamp 1626908933
transform 1 0 25152 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_904
timestamp 1626908933
transform 1 0 25152 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_905
timestamp 1626908933
transform 1 0 25152 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_246
timestamp 1626908933
transform 1 0 26400 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1237
timestamp 1626908933
transform 1 0 26400 0 -1 21312
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_56
timestamp 1626908933
transform 1 0 26900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_704
timestamp 1626908933
transform 1 0 26900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_56
timestamp 1626908933
transform 1 0 26900 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_704
timestamp 1626908933
transform 1 0 26900 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1252
timestamp 1626908933
transform 1 0 27264 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1236
timestamp 1626908933
transform 1 0 27264 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_261
timestamp 1626908933
transform 1 0 27264 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_245
timestamp 1626908933
transform 1 0 27264 0 -1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2313
timestamp 1626908933
transform 1 0 27312 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_378
timestamp 1626908933
transform 1 0 27312 0 1 19869
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1889
timestamp 1626908933
transform 1 0 27360 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_898
timestamp 1626908933
transform 1 0 27360 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_484
timestamp 1626908933
transform 1 0 27456 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_127
timestamp 1626908933
transform 1 0 27456 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_682
timestamp 1626908933
transform 1 0 27360 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_84
timestamp 1626908933
transform 1 0 27360 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_153
timestamp 1626908933
transform 1 0 26496 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_154
timestamp 1626908933
transform 1 0 26496 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_875
timestamp 1626908933
transform 1 0 26496 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_876
timestamp 1626908933
transform 1 0 26496 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_17
timestamp 1626908933
transform 1 0 27552 0 -1 21312
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_5
timestamp 1626908933
transform 1 0 27552 0 -1 21312
box -38 -49 1862 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1017
timestamp 1626908933
transform 1 0 28100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_369
timestamp 1626908933
transform 1 0 28100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1017
timestamp 1626908933
transform 1 0 28100 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_369
timestamp 1626908933
transform 1 0 28100 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_845
timestamp 1626908933
transform 1 0 27744 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_123
timestamp 1626908933
transform 1 0 27744 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_260
timestamp 1626908933
transform 1 0 28896 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1251
timestamp 1626908933
transform 1 0 28896 0 1 19980
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_32
timestamp 1626908933
transform 1 0 29300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_680
timestamp 1626908933
transform 1 0 29300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_32
timestamp 1626908933
transform 1 0 29300 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_680
timestamp 1626908933
transform 1 0 29300 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_88
timestamp 1626908933
transform 1 0 28992 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_810
timestamp 1626908933
transform 1 0 28992 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_60
timestamp 1626908933
transform 1 0 28512 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_658
timestamp 1626908933
transform 1 0 28512 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_131
timestamp 1626908933
transform 1 0 29376 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_732
timestamp 1626908933
transform 1 0 29376 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_259
timestamp 1626908933
transform 1 0 29760 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1250
timestamp 1626908933
transform 1 0 29760 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_133
timestamp 1626908933
transform 1 0 29952 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_490
timestamp 1626908933
transform 1 0 29952 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_136
timestamp 1626908933
transform 1 0 30048 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_737
timestamp 1626908933
transform 1 0 30048 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_891
timestamp 1626908933
transform 1 0 29856 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1882
timestamp 1626908933
transform 1 0 29856 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_73
timestamp 1626908933
transform 1 0 29568 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_795
timestamp 1626908933
transform 1 0 29568 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_27
timestamp 1626908933
transform 1 0 30336 0 -1 21312
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_12
timestamp 1626908933
transform 1 0 30336 0 -1 21312
box -38 -49 710 715
use L1M1_PR  L1M1_PR_2311
timestamp 1626908933
transform 1 0 30384 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_376
timestamp 1626908933
transform 1 0 30384 0 1 19869
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1249
timestamp 1626908933
transform 1 0 30240 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_258
timestamp 1626908933
transform 1 0 30240 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_764
timestamp 1626908933
transform 1 0 30336 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_42
timestamp 1626908933
transform 1 0 30336 0 1 19980
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_345
timestamp 1626908933
transform 1 0 30500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_993
timestamp 1626908933
transform 1 0 30500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_345
timestamp 1626908933
transform 1 0 30500 0 1 19980
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_993
timestamp 1626908933
transform 1 0 30500 0 1 19980
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_244
timestamp 1626908933
transform 1 0 31008 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_257
timestamp 1626908933
transform 1 0 31104 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1235
timestamp 1626908933
transform 1 0 31008 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1248
timestamp 1626908933
transform 1 0 31104 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_8
timestamp 1626908933
transform 1 0 31200 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_730
timestamp 1626908933
transform 1 0 31200 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_5
timestamp 1626908933
transform 1 0 31104 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_603
timestamp 1626908933
transform 1 0 31104 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_243
timestamp 1626908933
transform 1 0 31488 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1234
timestamp 1626908933
transform 1 0 31488 0 -1 21312
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_656
timestamp 1626908933
transform 1 0 31700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_8
timestamp 1626908933
transform 1 0 31700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_656
timestamp 1626908933
transform 1 0 31700 0 1 20646
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_8
timestamp 1626908933
transform 1 0 31700 0 1 20646
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1890
timestamp 1626908933
transform 1 0 31584 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_899
timestamp 1626908933
transform 1 0 31584 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1136
timestamp 1626908933
transform 1 0 31776 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_535
timestamp 1626908933
transform 1 0 31776 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_483
timestamp 1626908933
transform 1 0 31680 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_126
timestamp 1626908933
transform 1 0 31680 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_892
timestamp 1626908933
transform 1 0 31968 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_900
timestamp 1626908933
transform 1 0 31968 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1883
timestamp 1626908933
transform 1 0 31968 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1891
timestamp 1626908933
transform 1 0 31968 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_536
timestamp 1626908933
transform 1 0 0 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1137
timestamp 1626908933
transform 1 0 0 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_901
timestamp 1626908933
transform 1 0 192 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1892
timestamp 1626908933
transform 1 0 192 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_125
timestamp 1626908933
transform 1 0 288 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_482
timestamp 1626908933
transform 1 0 288 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_537
timestamp 1626908933
transform 1 0 384 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1138
timestamp 1626908933
transform 1 0 384 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_902
timestamp 1626908933
transform 1 0 576 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1893
timestamp 1626908933
transform 1 0 576 0 1 21312
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1280
timestamp 1626908933
transform 1 0 1700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_632
timestamp 1626908933
transform 1 0 1700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1280
timestamp 1626908933
transform 1 0 1700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_632
timestamp 1626908933
transform 1 0 1700 0 1 21312
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3099
timestamp 1626908933
transform 1 0 1584 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2947
timestamp 1626908933
transform 1 0 1392 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1132
timestamp 1626908933
transform 1 0 1584 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_980
timestamp 1626908933
transform 1 0 1392 0 1 20757
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_52
timestamp 1626908933
transform 1 0 672 0 1 21312
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_6
timestamp 1626908933
transform 1 0 672 0 1 21312
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_978
timestamp 1626908933
transform 1 0 3120 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2945
timestamp 1626908933
transform 1 0 3120 0 1 20757
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1041
timestamp 1626908933
transform 1 0 3120 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2976
timestamp 1626908933
transform 1 0 3120 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_302
timestamp 1626908933
transform 1 0 3312 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1129
timestamp 1626908933
transform 1 0 3120 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2269
timestamp 1626908933
transform 1 0 3312 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3096
timestamp 1626908933
transform 1 0 3120 0 1 21201
box -32 -32 32 32
use L1M1_PR  L1M1_PR_326
timestamp 1626908933
transform 1 0 3216 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1201
timestamp 1626908933
transform 1 0 3024 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2261
timestamp 1626908933
transform 1 0 3216 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3136
timestamp 1626908933
transform 1 0 3024 0 1 21053
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_641
timestamp 1626908933
transform 1 0 3360 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1363
timestamp 1626908933
transform 1 0 3360 0 1 21312
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2437
timestamp 1626908933
transform 1 0 4272 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_502
timestamp 1626908933
transform 1 0 4272 0 1 20905
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3838
timestamp 1626908933
transform 1 0 4176 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1871
timestamp 1626908933
transform 1 0 4176 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_472
timestamp 1626908933
transform 1 0 4272 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2439
timestamp 1626908933
transform 1 0 4272 0 1 21053
box -32 -32 32 32
use L1M1_PR  L1M1_PR_324
timestamp 1626908933
transform 1 0 4080 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2259
timestamp 1626908933
transform 1 0 4080 0 1 21053
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1859
timestamp 1626908933
transform 1 0 3984 0 1 21127
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3826
timestamp 1626908933
transform 1 0 3984 0 1 21127
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_608
timestamp 1626908933
transform 1 0 4100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1256
timestamp 1626908933
transform 1 0 4100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_608
timestamp 1626908933
transform 1 0 4100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1256
timestamp 1626908933
transform 1 0 4100 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1139
timestamp 1626908933
transform 1 0 4128 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_538
timestamp 1626908933
transform 1 0 4128 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_99
timestamp 1626908933
transform -1 0 4608 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_38
timestamp 1626908933
transform -1 0 4608 0 1 21312
box -38 -49 326 715
use L1M1_PR  L1M1_PR_468
timestamp 1626908933
transform 1 0 4368 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2403
timestamp 1626908933
transform 1 0 4368 0 1 21053
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1140
timestamp 1626908933
transform 1 0 5088 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_539
timestamp 1626908933
transform 1 0 5088 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1114
timestamp 1626908933
transform 1 0 4608 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_516
timestamp 1626908933
transform 1 0 4608 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_481
timestamp 1626908933
transform 1 0 4992 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_124
timestamp 1626908933
transform 1 0 4992 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_57
timestamp 1626908933
transform -1 0 5760 0 1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_126
timestamp 1626908933
transform -1 0 5760 0 1 21312
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3779
timestamp 1626908933
transform 1 0 5424 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3778
timestamp 1626908933
transform 1 0 5424 0 1 21201
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1844
timestamp 1626908933
transform 1 0 5424 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1843
timestamp 1626908933
transform 1 0 5424 0 1 21201
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3835
timestamp 1626908933
transform 1 0 5424 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1868
timestamp 1626908933
transform 1 0 5424 0 1 21201
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3769
timestamp 1626908933
transform 1 0 5712 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2439
timestamp 1626908933
transform 1 0 5616 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1834
timestamp 1626908933
transform 1 0 5712 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_504
timestamp 1626908933
transform 1 0 5616 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2475
timestamp 1626908933
transform 1 0 5616 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_508
timestamp 1626908933
transform 1 0 5616 0 1 20757
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_94
timestamp 1626908933
transform 1 0 5760 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_42
timestamp 1626908933
transform 1 0 5760 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_903
timestamp 1626908933
transform 1 0 6144 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1894
timestamp 1626908933
transform 1 0 6144 0 1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_506
timestamp 1626908933
transform 1 0 6288 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2473
timestamp 1626908933
transform 1 0 6288 0 1 20905
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2369
timestamp 1626908933
transform 1 0 6576 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_434
timestamp 1626908933
transform 1 0 6576 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2405
timestamp 1626908933
transform 1 0 6576 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_438
timestamp 1626908933
transform 1 0 6576 0 1 20757
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1232
timestamp 1626908933
transform 1 0 6500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_584
timestamp 1626908933
transform 1 0 6500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1232
timestamp 1626908933
transform 1 0 6500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_584
timestamp 1626908933
transform 1 0 6500 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1233
timestamp 1626908933
transform 1 0 6528 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_242
timestamp 1626908933
transform 1 0 6528 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_480
timestamp 1626908933
transform 1 0 6624 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1078
timestamp 1626908933
transform 1 0 6624 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_0
timestamp 1626908933
transform 1 0 6240 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_62
timestamp 1626908933
transform 1 0 6240 0 1 21312
box -38 -49 326 715
use M1M2_PR  M1M2_PR_2416
timestamp 1626908933
transform 1 0 6960 0 1 20831
box -32 -32 32 32
use M1M2_PR  M1M2_PR_449
timestamp 1626908933
transform 1 0 6960 0 1 20831
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3762
timestamp 1626908933
transform 1 0 6864 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1827
timestamp 1626908933
transform 1 0 6864 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3817
timestamp 1626908933
transform 1 0 6768 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1850
timestamp 1626908933
transform 1 0 6768 0 1 20979
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2371
timestamp 1626908933
transform 1 0 6960 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_436
timestamp 1626908933
transform 1 0 6960 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2408
timestamp 1626908933
transform 1 0 6960 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_441
timestamp 1626908933
transform 1 0 6960 0 1 20979
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2373
timestamp 1626908933
transform 1 0 7152 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_438
timestamp 1626908933
transform 1 0 7152 0 1 20905
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2409
timestamp 1626908933
transform 1 0 7152 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_442
timestamp 1626908933
transform 1 0 7152 0 1 20905
box -32 -32 32 32
use L1M1_PR  L1M1_PR_433
timestamp 1626908933
transform 1 0 6960 0 1 21201
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2368
timestamp 1626908933
transform 1 0 6960 0 1 21201
box -29 -23 29 23
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_0
timestamp 1626908933
transform 1 0 7008 0 1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__o21ai_1  sky130_fd_sc_hs__o21ai_1_6
timestamp 1626908933
transform 1 0 7008 0 1 21312
box -38 -49 518 715
use M1M2_PR  M1M2_PR_2404
timestamp 1626908933
transform 1 0 7344 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2251
timestamp 1626908933
transform 1 0 7344 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_437
timestamp 1626908933
transform 1 0 7344 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_284
timestamp 1626908933
transform 1 0 7344 0 1 20979
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_95
timestamp 1626908933
transform 1 0 7488 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_43
timestamp 1626908933
transform 1 0 7488 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1895
timestamp 1626908933
transform 1 0 7872 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_904
timestamp 1626908933
transform 1 0 7872 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_56
timestamp 1626908933
transform 1 0 7968 0 1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_125
timestamp 1626908933
transform 1 0 7968 0 1 21312
box -38 -49 518 715
use M1M2_PR  M1M2_PR_3169
timestamp 1626908933
transform 1 0 8304 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1202
timestamp 1626908933
transform 1 0 8304 0 1 20757
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3205
timestamp 1626908933
transform 1 0 8592 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1270
timestamp 1626908933
transform 1 0 8592 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2397
timestamp 1626908933
transform 1 0 9072 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_462
timestamp 1626908933
transform 1 0 9072 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2428
timestamp 1626908933
transform 1 0 9072 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_461
timestamp 1626908933
transform 1 0 9072 0 1 20757
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2241
timestamp 1626908933
transform 1 0 8400 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_306
timestamp 1626908933
transform 1 0 8400 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2249
timestamp 1626908933
transform 1 0 8688 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_282
timestamp 1626908933
transform 1 0 8688 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_455
timestamp 1626908933
transform 1 0 8496 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2422
timestamp 1626908933
transform 1 0 8496 0 1 21053
box -32 -32 32 32
use L1M1_PR  L1M1_PR_456
timestamp 1626908933
transform 1 0 8304 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2391
timestamp 1626908933
transform 1 0 8304 0 1 21053
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_560
timestamp 1626908933
transform 1 0 8900 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1208
timestamp 1626908933
transform 1 0 8900 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_560
timestamp 1626908933
transform 1 0 8900 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1208
timestamp 1626908933
transform 1 0 8900 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_548
timestamp 1626908933
transform 1 0 8448 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1270
timestamp 1626908933
transform 1 0 8448 0 1 21312
box -38 -49 806 715
use M1M2_PR  M1M2_PR_225
timestamp 1626908933
transform 1 0 9552 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2192
timestamp 1626908933
transform 1 0 9552 0 1 20757
box -32 -32 32 32
use L1M1_PR  L1M1_PR_449
timestamp 1626908933
transform 1 0 9456 0 1 20831
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2384
timestamp 1626908933
transform 1 0 9456 0 1 20831
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_123
timestamp 1626908933
transform 1 0 9984 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_480
timestamp 1626908933
transform 1 0 9984 0 1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_198
timestamp 1626908933
transform 1 0 9648 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2165
timestamp 1626908933
transform 1 0 9648 0 1 20979
box -32 -32 32 32
use L1M1_PR  L1M1_PR_217
timestamp 1626908933
transform 1 0 9648 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_453
timestamp 1626908933
transform 1 0 9744 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2152
timestamp 1626908933
transform 1 0 9648 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2388
timestamp 1626908933
transform 1 0 9744 0 1 21053
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_525
timestamp 1626908933
transform 1 0 9216 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1247
timestamp 1626908933
transform 1 0 9216 0 1 21312
box -38 -49 806 715
use L1M1_PR  L1M1_PR_245
timestamp 1626908933
transform 1 0 10320 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2180
timestamp 1626908933
transform 1 0 10320 0 1 20757
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_241
timestamp 1626908933
transform 1 0 10656 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1232
timestamp 1626908933
transform 1 0 10656 0 1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1090
timestamp 1626908933
transform 1 0 10800 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3025
timestamp 1626908933
transform 1 0 10800 0 1 20979
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_493
timestamp 1626908933
transform 1 0 10752 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1215
timestamp 1626908933
transform 1 0 10752 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_5
timestamp 1626908933
transform 1 0 10080 0 1 21312
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_18
timestamp 1626908933
transform 1 0 10080 0 1 21312
box -38 -49 614 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_536
timestamp 1626908933
transform 1 0 11300 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1184
timestamp 1626908933
transform 1 0 11300 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_536
timestamp 1626908933
transform 1 0 11300 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1184
timestamp 1626908933
transform 1 0 11300 0 1 21312
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3604
timestamp 1626908933
transform 1 0 11760 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1669
timestamp 1626908933
transform 1 0 11760 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3547
timestamp 1626908933
transform 1 0 11472 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2990
timestamp 1626908933
transform 1 0 11472 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1580
timestamp 1626908933
transform 1 0 11472 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1023
timestamp 1626908933
transform 1 0 11472 0 1 20979
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3029
timestamp 1626908933
transform 1 0 11664 0 1 21201
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1094
timestamp 1626908933
transform 1 0 11664 0 1 21201
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_112
timestamp 1626908933
transform 1 0 11520 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_50
timestamp 1626908933
transform 1 0 11520 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_130
timestamp 1626908933
transform 1 0 11808 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_731
timestamp 1626908933
transform 1 0 11808 0 1 21312
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1027
timestamp 1626908933
transform 1 0 11856 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2994
timestamp 1626908933
transform 1 0 11856 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1564
timestamp 1626908933
transform 1 0 12144 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3531
timestamp 1626908933
transform 1 0 12144 0 1 20757
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1088
timestamp 1626908933
transform 1 0 11952 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3023
timestamp 1626908933
transform 1 0 11952 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1020
timestamp 1626908933
transform 1 0 12048 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2987
timestamp 1626908933
transform 1 0 12048 0 1 21053
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1085
timestamp 1626908933
transform 1 0 12048 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3020
timestamp 1626908933
transform 1 0 12048 0 1 21053
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_470
timestamp 1626908933
transform 1 0 12000 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1192
timestamp 1626908933
transform 1 0 12000 0 1 21312
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3588
timestamp 1626908933
transform 1 0 13008 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1653
timestamp 1626908933
transform 1 0 13008 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3033
timestamp 1626908933
transform 1 0 12912 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1066
timestamp 1626908933
transform 1 0 12912 0 1 20979
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3072
timestamp 1626908933
transform 1 0 13008 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1137
timestamp 1626908933
transform 1 0 13008 0 1 21053
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3038
timestamp 1626908933
transform 1 0 13008 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3032
timestamp 1626908933
transform 1 0 13104 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1071
timestamp 1626908933
transform 1 0 13008 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1065
timestamp 1626908933
transform 1 0 13104 0 1 21053
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_108
timestamp 1626908933
transform 1 0 12768 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_46
timestamp 1626908933
transform 1 0 12768 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_730
timestamp 1626908933
transform 1 0 13056 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_129
timestamp 1626908933
transform 1 0 13056 0 1 21312
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1130
timestamp 1626908933
transform 1 0 13296 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1133
timestamp 1626908933
transform 1 0 13200 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3065
timestamp 1626908933
transform 1 0 13296 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3068
timestamp 1626908933
transform 1 0 13200 0 1 20979
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_439
timestamp 1626908933
transform 1 0 13248 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1161
timestamp 1626908933
transform 1 0 13248 0 1 21312
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1160
timestamp 1626908933
transform 1 0 13700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_512
timestamp 1626908933
transform 1 0 13700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1160
timestamp 1626908933
transform 1 0 13700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_512
timestamp 1626908933
transform 1 0 13700 0 1 21312
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2211
timestamp 1626908933
transform 1 0 14640 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_276
timestamp 1626908933
transform 1 0 14640 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2220
timestamp 1626908933
transform 1 0 14640 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_253
timestamp 1626908933
transform 1 0 14640 0 1 20979
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_96
timestamp 1626908933
transform 1 0 14304 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_44
timestamp 1626908933
transform 1 0 14304 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_107
timestamp 1626908933
transform 1 0 14016 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_46
timestamp 1626908933
transform 1 0 14016 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_122
timestamp 1626908933
transform 1 0 14976 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_479
timestamp 1626908933
transform 1 0 14976 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_540
timestamp 1626908933
transform 1 0 14688 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1141
timestamp 1626908933
transform 1 0 14688 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_905
timestamp 1626908933
transform 1 0 14880 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1896
timestamp 1626908933
transform 1 0 14880 0 1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1132
timestamp 1626908933
transform 1 0 14736 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3067
timestamp 1626908933
transform 1 0 14736 0 1 20905
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_240
timestamp 1626908933
transform 1 0 15456 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1231
timestamp 1626908933
transform 1 0 15456 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_316
timestamp 1626908933
transform 1 0 15072 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_914
timestamp 1626908933
transform 1 0 15072 0 1 21312
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1136
timestamp 1626908933
transform 1 0 16100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_488
timestamp 1626908933
transform 1 0 16100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1136
timestamp 1626908933
transform 1 0 16100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_488
timestamp 1626908933
transform 1 0 16100 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1230
timestamp 1626908933
transform 1 0 16320 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_239
timestamp 1626908933
transform 1 0 16320 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1127
timestamp 1626908933
transform 1 0 15552 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_405
timestamp 1626908933
transform 1 0 15552 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_69
timestamp 1626908933
transform -1 0 17088 0 1 21312
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_30
timestamp 1626908933
transform -1 0 17088 0 1 21312
box -38 -49 614 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1897
timestamp 1626908933
transform 1 0 16416 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_906
timestamp 1626908933
transform 1 0 16416 0 1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1979
timestamp 1626908933
transform 1 0 17520 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_12
timestamp 1626908933
transform 1 0 17520 0 1 20979
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_729
timestamp 1626908933
transform 1 0 17088 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_128
timestamp 1626908933
transform 1 0 17088 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1089
timestamp 1626908933
transform 1 0 17280 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_367
timestamp 1626908933
transform 1 0 17280 0 1 21312
box -38 -49 806 715
use L1M1_PR  L1M1_PR_14
timestamp 1626908933
transform 1 0 18000 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1949
timestamp 1626908933
transform 1 0 18000 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1536
timestamp 1626908933
transform 1 0 18192 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3503
timestamp 1626908933
transform 1 0 18192 0 1 21053
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1623
timestamp 1626908933
transform 1 0 18192 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3558
timestamp 1626908933
transform 1 0 18192 0 1 21053
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_464
timestamp 1626908933
transform 1 0 18500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1112
timestamp 1626908933
transform 1 0 18500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_464
timestamp 1626908933
transform 1 0 18500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1112
timestamp 1626908933
transform 1 0 18500 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_133
timestamp 1626908933
transform -1 0 18528 0 1 21312
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_64
timestamp 1626908933
transform -1 0 18528 0 1 21312
box -38 -49 518 715
use M1M2_PR  M1M2_PR_2362
timestamp 1626908933
transform 1 0 19056 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_395
timestamp 1626908933
transform 1 0 19056 0 1 20905
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1898
timestamp 1626908933
transform 1 0 18720 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_907
timestamp 1626908933
transform 1 0 18720 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1142
timestamp 1626908933
transform 1 0 18528 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_541
timestamp 1626908933
transform 1 0 18528 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__nor2_4  sky130_fd_sc_hs__nor2_4_2
timestamp 1626908933
transform -1 0 19680 0 1 21312
box -38 -49 902 715
use sky130_fd_sc_hs__nor2_4  sky130_fd_sc_hs__nor2_4_0
timestamp 1626908933
transform -1 0 19680 0 1 21312
box -38 -49 902 715
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_2
timestamp 1626908933
transform 1 0 19680 0 1 21312
box -38 -49 326 715
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_0
timestamp 1626908933
transform 1 0 19680 0 1 21312
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1433
timestamp 1626908933
transform 1 0 19632 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3400
timestamp 1626908933
transform 1 0 19632 0 1 20905
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_121
timestamp 1626908933
transform 1 0 19968 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_478
timestamp 1626908933
transform 1 0 19968 0 1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1517
timestamp 1626908933
transform 1 0 20016 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3452
timestamp 1626908933
transform 1 0 20016 0 1 20905
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1313
timestamp 1626908933
transform 1 0 20112 0 1 21127
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1395
timestamp 1626908933
transform 1 0 20304 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3280
timestamp 1626908933
transform 1 0 20112 0 1 21127
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3362
timestamp 1626908933
transform 1 0 20304 0 1 21201
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1088
timestamp 1626908933
transform 1 0 20900 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_440
timestamp 1626908933
transform 1 0 20900 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1088
timestamp 1626908933
transform 1 0 20900 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_440
timestamp 1626908933
transform 1 0 20900 0 1 21312
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3327
timestamp 1626908933
transform 1 0 21360 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1392
timestamp 1626908933
transform 1 0 21360 0 1 21053
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3396
timestamp 1626908933
transform 1 0 21456 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1429
timestamp 1626908933
transform 1 0 21456 0 1 21053
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3449
timestamp 1626908933
transform 1 0 21552 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3412
timestamp 1626908933
transform 1 0 21552 0 1 21201
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1514
timestamp 1626908933
transform 1 0 21552 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1477
timestamp 1626908933
transform 1 0 21552 0 1 21201
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_269
timestamp 1626908933
transform 1 0 21984 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_991
timestamp 1626908933
transform 1 0 21984 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__sdlclkp_4  sky130_fd_sc_hs__sdlclkp_4_1
timestamp 1626908933
transform 1 0 20064 0 1 21312
box -38 -49 1958 715
use sky130_fd_sc_hs__sdlclkp_4  sky130_fd_sc_hs__sdlclkp_4_0
timestamp 1626908933
transform 1 0 20064 0 1 21312
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_2301
timestamp 1626908933
transform 1 0 22608 0 1 21201
box -32 -32 32 32
use M1M2_PR  M1M2_PR_334
timestamp 1626908933
transform 1 0 22608 0 1 21201
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_768
timestamp 1626908933
transform 1 0 22752 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_170
timestamp 1626908933
transform 1 0 22752 0 1 21312
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3357
timestamp 1626908933
transform 1 0 23088 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1422
timestamp 1626908933
transform 1 0 23088 0 1 20757
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3307
timestamp 1626908933
transform 1 0 23088 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1340
timestamp 1626908933
transform 1 0 23088 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3237
timestamp 1626908933
transform 1 0 23088 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1270
timestamp 1626908933
transform 1 0 23088 0 1 20905
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3291
timestamp 1626908933
transform 1 0 23280 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1356
timestamp 1626908933
transform 1 0 23280 0 1 20905
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1064
timestamp 1626908933
transform 1 0 23300 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_416
timestamp 1626908933
transform 1 0 23300 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1064
timestamp 1626908933
transform 1 0 23300 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_416
timestamp 1626908933
transform 1 0 23300 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_238
timestamp 1626908933
transform 1 0 23808 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1229
timestamp 1626908933
transform 1 0 23808 0 1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1303
timestamp 1626908933
transform 1 0 23472 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1426
timestamp 1626908933
transform 1 0 23664 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3270
timestamp 1626908933
transform 1 0 23472 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3393
timestamp 1626908933
transform 1 0 23664 0 1 21053
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_1
timestamp 1626908933
transform 1 0 23136 0 1 21312
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_16
timestamp 1626908933
transform 1 0 23136 0 1 21312
box -38 -49 710 715
use M1M2_PR  M1M2_PR_370
timestamp 1626908933
transform 1 0 24144 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1271
timestamp 1626908933
transform 1 0 24048 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2337
timestamp 1626908933
transform 1 0 24144 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3238
timestamp 1626908933
transform 1 0 24048 0 1 20905
box -32 -32 32 32
use L1M1_PR  L1M1_PR_392
timestamp 1626908933
transform 1 0 24624 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1358
timestamp 1626908933
transform 1 0 24048 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2327
timestamp 1626908933
transform 1 0 24624 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3293
timestamp 1626908933
transform 1 0 24048 0 1 20905
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_216
timestamp 1626908933
transform 1 0 23904 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_938
timestamp 1626908933
transform 1 0 23904 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1228
timestamp 1626908933
transform 1 0 24864 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_237
timestamp 1626908933
transform 1 0 24864 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_728
timestamp 1626908933
transform 1 0 24672 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_127
timestamp 1626908933
transform 1 0 24672 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_120
timestamp 1626908933
transform 1 0 24960 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_477
timestamp 1626908933
transform 1 0 24960 0 1 21312
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_392
timestamp 1626908933
transform 1 0 25700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1040
timestamp 1626908933
transform 1 0 25700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_392
timestamp 1626908933
transform 1 0 25700 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1040
timestamp 1626908933
transform 1 0 25700 0 1 21312
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1406
timestamp 1626908933
transform 1 0 25872 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1424
timestamp 1626908933
transform 1 0 25872 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3373
timestamp 1626908933
transform 1 0 25872 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3391
timestamp 1626908933
transform 1 0 25872 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1278
timestamp 1626908933
transform 1 0 26064 0 1 20831
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3245
timestamp 1626908933
transform 1 0 26064 0 1 20831
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1489
timestamp 1626908933
transform 1 0 25968 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3424
timestamp 1626908933
transform 1 0 25968 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1508
timestamp 1626908933
transform 1 0 26160 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3443
timestamp 1626908933
transform 1 0 26160 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3367
timestamp 1626908933
transform 1 0 26352 0 1 21053
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1432
timestamp 1626908933
transform 1 0 26352 0 1 21053
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3267
timestamp 1626908933
transform 1 0 26736 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1300
timestamp 1626908933
transform 1 0 26736 0 1 20979
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_48
timestamp 1626908933
transform 1 0 25056 0 1 21312
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_2
timestamp 1626908933
transform 1 0 25056 0 1 21312
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_353
timestamp 1626908933
transform 1 0 27696 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1295
timestamp 1626908933
transform 1 0 28464 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2320
timestamp 1626908933
transform 1 0 27696 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3262
timestamp 1626908933
transform 1 0 28464 0 1 20979
box -32 -32 32 32
use L1M1_PR  L1M1_PR_377
timestamp 1626908933
transform 1 0 27696 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1368
timestamp 1626908933
transform 1 0 27984 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2312
timestamp 1626908933
transform 1 0 27696 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3303
timestamp 1626908933
transform 1 0 27984 0 1 20905
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_368
timestamp 1626908933
transform 1 0 28100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1016
timestamp 1626908933
transform 1 0 28100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_368
timestamp 1626908933
transform 1 0 28100 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1016
timestamp 1626908933
transform 1 0 28100 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_122
timestamp 1626908933
transform 1 0 27744 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_844
timestamp 1626908933
transform 1 0 27744 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_908
timestamp 1626908933
transform 1 0 28512 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1899
timestamp 1626908933
transform 1 0 28512 0 1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3301
timestamp 1626908933
transform 1 0 29040 0 1 20905
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1366
timestamp 1626908933
transform 1 0 29040 0 1 20905
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3242
timestamp 1626908933
transform 1 0 28944 0 1 20905
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1275
timestamp 1626908933
transform 1 0 28944 0 1 20905
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3366
timestamp 1626908933
transform 1 0 29232 0 1 21127
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1431
timestamp 1626908933
transform 1 0 29232 0 1 21127
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3858
timestamp 1626908933
transform 1 0 29040 0 1 21053
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1891
timestamp 1626908933
transform 1 0 29040 0 1 21053
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_727
timestamp 1626908933
transform 1 0 29280 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_126
timestamp 1626908933
transform 1 0 29280 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_7
timestamp 1626908933
transform 1 0 28608 0 1 21312
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_22
timestamp 1626908933
transform 1 0 28608 0 1 21312
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1227
timestamp 1626908933
transform 1 0 29472 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_236
timestamp 1626908933
transform 1 0 29472 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_726
timestamp 1626908933
transform 1 0 30048 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_125
timestamp 1626908933
transform 1 0 30048 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_639
timestamp 1626908933
transform 1 0 29568 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_41
timestamp 1626908933
transform 1 0 29568 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_476
timestamp 1626908933
transform 1 0 29952 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_119
timestamp 1626908933
transform 1 0 29952 0 1 21312
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3744
timestamp 1626908933
transform 1 0 30288 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2294
timestamp 1626908933
transform 1 0 30384 0 1 21201
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1809
timestamp 1626908933
transform 1 0 30288 0 1 20757
box -29 -23 29 23
use L1M1_PR  L1M1_PR_359
timestamp 1626908933
transform 1 0 30384 0 1 21201
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1226
timestamp 1626908933
transform 1 0 30240 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_235
timestamp 1626908933
transform 1 0 30240 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_763
timestamp 1626908933
transform 1 0 30336 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_41
timestamp 1626908933
transform 1 0 30336 0 1 21312
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3791
timestamp 1626908933
transform 1 0 30768 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2338
timestamp 1626908933
transform 1 0 30672 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1856
timestamp 1626908933
transform 1 0 30768 0 1 20979
box -29 -23 29 23
use L1M1_PR  L1M1_PR_403
timestamp 1626908933
transform 1 0 30672 0 1 20979
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3848
timestamp 1626908933
transform 1 0 30768 0 1 20831
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2377
timestamp 1626908933
transform 1 0 30672 0 1 20979
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1881
timestamp 1626908933
transform 1 0 30768 0 1 20831
box -32 -32 32 32
use M1M2_PR  M1M2_PR_410
timestamp 1626908933
transform 1 0 30672 0 1 20979
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_992
timestamp 1626908933
transform 1 0 30500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_344
timestamp 1626908933
transform 1 0 30500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_992
timestamp 1626908933
transform 1 0 30500 0 1 21312
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_344
timestamp 1626908933
transform 1 0 30500 0 1 21312
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_234
timestamp 1626908933
transform 1 0 31104 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1225
timestamp 1626908933
transform 1 0 31104 0 1 21312
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1773
timestamp 1626908933
transform 1 0 31152 0 1 20831
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3740
timestamp 1626908933
transform 1 0 31152 0 1 20831
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1790
timestamp 1626908933
transform 1 0 30960 0 1 20831
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3725
timestamp 1626908933
transform 1 0 30960 0 1 20831
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_7
timestamp 1626908933
transform 1 0 31200 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_729
timestamp 1626908933
transform 1 0 31200 0 1 21312
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3781
timestamp 1626908933
transform 1 0 31920 0 1 20757
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1814
timestamp 1626908933
transform 1 0 31920 0 1 20757
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1900
timestamp 1626908933
transform 1 0 31968 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_909
timestamp 1626908933
transform 1 0 31968 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_124
timestamp 1626908933
transform 1 0 0 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_725
timestamp 1626908933
transform 1 0 0 0 -1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1854
timestamp 1626908933
transform 1 0 48 0 1 21793
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3821
timestamp 1626908933
transform 1 0 48 0 1 21793
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1628
timestamp 1626908933
transform 1 0 720 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3563
timestamp 1626908933
transform 1 0 720 0 1 21571
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_319
timestamp 1626908933
transform 1 0 500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_967
timestamp 1626908933
transform 1 0 500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_319
timestamp 1626908933
transform 1 0 500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_967
timestamp 1626908933
transform 1 0 500 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_707
timestamp 1626908933
transform 1 0 192 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1429
timestamp 1626908933
transform 1 0 192 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_233
timestamp 1626908933
transform 1 0 960 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1224
timestamp 1626908933
transform 1 0 960 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1540
timestamp 1626908933
transform 1 0 1200 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3507
timestamp 1626908933
transform 1 0 1200 0 1 21571
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1730
timestamp 1626908933
transform 1 0 1104 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3665
timestamp 1626908933
transform 1 0 1104 0 1 21645
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_673
timestamp 1626908933
transform 1 0 1440 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1395
timestamp 1626908933
transform 1 0 1440 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_569
timestamp 1626908933
transform 1 0 1056 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1167
timestamp 1626908933
transform 1 0 1056 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_232
timestamp 1626908933
transform 1 0 2208 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1223
timestamp 1626908933
transform 1 0 2208 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1173
timestamp 1626908933
transform 1 0 2064 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3140
timestamp 1626908933
transform 1 0 2064 0 1 21719
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_118
timestamp 1626908933
transform 1 0 2496 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_475
timestamp 1626908933
transform 1 0 2496 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_542
timestamp 1626908933
transform 1 0 2304 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1143
timestamp 1626908933
transform 1 0 2304 0 -1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1172
timestamp 1626908933
transform 1 0 2448 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3139
timestamp 1626908933
transform 1 0 2448 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3612
timestamp 1626908933
transform 1 0 2736 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1645
timestamp 1626908933
transform 1 0 2736 0 1 21645
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_97
timestamp 1626908933
transform 1 0 2592 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_45
timestamp 1626908933
transform 1 0 2592 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_910
timestamp 1626908933
transform 1 0 2976 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1901
timestamp 1626908933
transform 1 0 2976 0 -1 22644
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_295
timestamp 1626908933
transform 1 0 2900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_943
timestamp 1626908933
transform 1 0 2900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_295
timestamp 1626908933
transform 1 0 2900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_943
timestamp 1626908933
transform 1 0 2900 0 1 21978
box -100 -49 100 49
use M1M2_PR  M1M2_PR_301
timestamp 1626908933
transform 1 0 3312 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1115
timestamp 1626908933
transform 1 0 3312 0 1 21793
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2268
timestamp 1626908933
transform 1 0 3312 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3082
timestamp 1626908933
transform 1 0 3312 0 1 21793
box -32 -32 32 32
use L1M1_PR  L1M1_PR_325
timestamp 1626908933
transform 1 0 3216 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1180
timestamp 1626908933
transform 1 0 3216 0 1 22089
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2260
timestamp 1626908933
transform 1 0 3216 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3115
timestamp 1626908933
transform 1 0 3216 0 1 22089
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_36
timestamp 1626908933
transform -1 0 3648 0 -1 22644
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_75
timestamp 1626908933
transform -1 0 3648 0 -1 22644
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2246
timestamp 1626908933
transform 1 0 4368 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_311
timestamp 1626908933
transform 1 0 4368 0 1 21571
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1124
timestamp 1626908933
transform 1 0 3648 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_526
timestamp 1626908933
transform 1 0 3648 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1349
timestamp 1626908933
transform 1 0 4032 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_627
timestamp 1626908933
transform 1 0 4032 0 -1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_289
timestamp 1626908933
transform 1 0 4464 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1110
timestamp 1626908933
transform 1 0 4560 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2256
timestamp 1626908933
transform 1 0 4464 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3077
timestamp 1626908933
transform 1 0 4560 0 1 21571
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1178
timestamp 1626908933
transform 1 0 4560 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3113
timestamp 1626908933
transform 1 0 4560 0 1 21571
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1109
timestamp 1626908933
transform 1 0 4560 0 1 22089
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3076
timestamp 1626908933
transform 1 0 4560 0 1 22089
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1182
timestamp 1626908933
transform 1 0 4464 0 1 21793
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3117
timestamp 1626908933
transform 1 0 4464 0 1 21793
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_271
timestamp 1626908933
transform 1 0 5300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_919
timestamp 1626908933
transform 1 0 5300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_271
timestamp 1626908933
transform 1 0 5300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_919
timestamp 1626908933
transform 1 0 5300 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_601
timestamp 1626908933
transform 1 0 4800 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1323
timestamp 1626908933
transform 1 0 4800 0 -1 22644
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3777
timestamp 1626908933
transform 1 0 5424 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1842
timestamp 1626908933
transform 1 0 5424 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3834
timestamp 1626908933
transform 1 0 5424 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1867
timestamp 1626908933
transform 1 0 5424 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1183
timestamp 1626908933
transform 1 0 5808 0 1 22163
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3150
timestamp 1626908933
transform 1 0 5808 0 1 22163
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1247
timestamp 1626908933
transform 1 0 5616 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1841
timestamp 1626908933
transform 1 0 5808 0 1 21719
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3182
timestamp 1626908933
transform 1 0 5616 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3776
timestamp 1626908933
transform 1 0 5808 0 1 21719
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3767
timestamp 1626908933
transform 1 0 6288 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1832
timestamp 1626908933
transform 1 0 6288 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3825
timestamp 1626908933
transform 1 0 6000 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1858
timestamp 1626908933
transform 1 0 6000 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3152
timestamp 1626908933
transform 1 0 6096 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2472
timestamp 1626908933
transform 1 0 6288 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1185
timestamp 1626908933
transform 1 0 6096 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_505
timestamp 1626908933
transform 1 0 6288 0 1 21867
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_724
timestamp 1626908933
transform 1 0 6240 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_123
timestamp 1626908933
transform 1 0 6240 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_4
timestamp 1626908933
transform 1 0 5568 0 -1 22644
box -38 -49 710 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_9
timestamp 1626908933
transform 1 0 5568 0 -1 22644
box -38 -49 710 715
use L1M1_PR  L1M1_PR_3774
timestamp 1626908933
transform 1 0 6480 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2372
timestamp 1626908933
transform 1 0 6384 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1839
timestamp 1626908933
transform 1 0 6480 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_437
timestamp 1626908933
transform 1 0 6384 0 1 21423
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1222
timestamp 1626908933
transform 1 0 6432 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_231
timestamp 1626908933
transform 1 0 6432 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3832
timestamp 1626908933
transform 1 0 6768 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3816
timestamp 1626908933
transform 1 0 6768 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1865
timestamp 1626908933
transform 1 0 6768 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1849
timestamp 1626908933
transform 1 0 6768 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_435
timestamp 1626908933
transform 1 0 7152 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_440
timestamp 1626908933
transform 1 0 6960 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2402
timestamp 1626908933
transform 1 0 7152 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2407
timestamp 1626908933
transform 1 0 6960 0 1 21423
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1826
timestamp 1626908933
transform 1 0 7056 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3761
timestamp 1626908933
transform 1 0 7056 0 1 21571
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_573
timestamp 1626908933
transform 1 0 6528 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1295
timestamp 1626908933
transform 1 0 6528 0 -1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_436
timestamp 1626908933
transform 1 0 7344 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2403
timestamp 1626908933
transform 1 0 7344 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_430
timestamp 1626908933
transform 1 0 7248 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_432
timestamp 1626908933
transform 1 0 7344 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2365
timestamp 1626908933
transform 1 0 7248 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2367
timestamp 1626908933
transform 1 0 7344 0 1 21645
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_230
timestamp 1626908933
transform 1 0 7296 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_911
timestamp 1626908933
transform 1 0 7392 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1221
timestamp 1626908933
transform 1 0 7296 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1902
timestamp 1626908933
transform 1 0 7392 0 -1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3559
timestamp 1626908933
transform 1 0 7440 0 1 21497
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1624
timestamp 1626908933
transform 1 0 7440 0 1 21497
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_474
timestamp 1626908933
transform 1 0 7488 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_117
timestamp 1626908933
transform 1 0 7488 0 -1 22644
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_895
timestamp 1626908933
transform 1 0 7700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_247
timestamp 1626908933
transform 1 0 7700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_895
timestamp 1626908933
transform 1 0 7700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_247
timestamp 1626908933
transform 1 0 7700 0 1 21978
box -100 -49 100 49
use L1M1_PR  L1M1_PR_500
timestamp 1626908933
transform 1 0 7920 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2435
timestamp 1626908933
transform 1 0 7920 0 1 21867
box -29 -23 29 23
use sky130_fd_sc_hs__a211oi_1  sky130_fd_sc_hs__a211oi_1_1
timestamp 1626908933
transform -1 0 8160 0 -1 22644
box -38 -49 614 715
use sky130_fd_sc_hs__a211oi_1  sky130_fd_sc_hs__a211oi_1_3
timestamp 1626908933
transform -1 0 8160 0 -1 22644
box -38 -49 614 715
use L1M1_PR  L1M1_PR_3195
timestamp 1626908933
transform 1 0 8112 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1260
timestamp 1626908933
transform 1 0 8112 0 1 21867
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3166
timestamp 1626908933
transform 1 0 8112 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1199
timestamp 1626908933
transform 1 0 8112 0 1 21867
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_40
timestamp 1626908933
transform 1 0 8160 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_17
timestamp 1626908933
transform 1 0 8160 0 -1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_454
timestamp 1626908933
transform 1 0 8496 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2421
timestamp 1626908933
transform 1 0 8496 0 1 21645
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_40
timestamp 1626908933
transform -1 0 9312 0 -1 22644
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_101
timestamp 1626908933
transform -1 0 9312 0 -1 22644
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_912
timestamp 1626908933
transform 1 0 8928 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1903
timestamp 1626908933
transform 1 0 8928 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_434
timestamp 1626908933
transform 1 0 9408 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1032
timestamp 1626908933
transform 1 0 9408 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_229
timestamp 1626908933
transform 1 0 9312 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1220
timestamp 1626908933
transform 1 0 9312 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1187
timestamp 1626908933
transform 1 0 9456 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3154
timestamp 1626908933
transform 1 0 9456 0 1 21719
box -32 -32 32 32
use L1M1_PR  L1M1_PR_452
timestamp 1626908933
transform 1 0 10128 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1248
timestamp 1626908933
transform 1 0 10224 0 1 21719
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2387
timestamp 1626908933
transform 1 0 10128 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3183
timestamp 1626908933
transform 1 0 10224 0 1 21719
box -29 -23 29 23
use M1M2_PR  M1M2_PR_217
timestamp 1626908933
transform 1 0 10320 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2184
timestamp 1626908933
transform 1 0 10320 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_235
timestamp 1626908933
transform 1 0 10320 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_267
timestamp 1626908933
transform 1 0 10416 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2170
timestamp 1626908933
transform 1 0 10320 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2202
timestamp 1626908933
transform 1 0 10416 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_489
timestamp 1626908933
transform 1 0 10512 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2456
timestamp 1626908933
transform 1 0 10512 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_486
timestamp 1626908933
transform 1 0 10512 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2421
timestamp 1626908933
transform 1 0 10512 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_488
timestamp 1626908933
transform 1 0 10896 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2455
timestamp 1626908933
transform 1 0 10896 0 1 21645
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_223
timestamp 1626908933
transform 1 0 10100 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_871
timestamp 1626908933
transform 1 0 10100 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_223
timestamp 1626908933
transform 1 0 10100 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_871
timestamp 1626908933
transform 1 0 10100 0 1 21978
box -100 -49 100 49
use L1M1_PR  L1M1_PR_236
timestamp 1626908933
transform 1 0 10224 0 1 22089
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2171
timestamp 1626908933
transform 1 0 10224 0 1 22089
box -29 -23 29 23
use M1M2_PR  M1M2_PR_216
timestamp 1626908933
transform 1 0 10320 0 1 22089
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2183
timestamp 1626908933
transform 1 0 10320 0 1 22089
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_75
timestamp 1626908933
transform -1 0 12480 0 -1 22644
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_29
timestamp 1626908933
transform -1 0 12480 0 -1 22644
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1022
timestamp 1626908933
transform 1 0 11472 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2989
timestamp 1626908933
transform 1 0 11472 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1086
timestamp 1626908933
transform 1 0 11760 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1089
timestamp 1626908933
transform 1 0 11568 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1093
timestamp 1626908933
transform 1 0 11664 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3021
timestamp 1626908933
transform 1 0 11760 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3024
timestamp 1626908933
transform 1 0 11568 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3028
timestamp 1626908933
transform 1 0 11664 0 1 21423
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1026
timestamp 1626908933
transform 1 0 11856 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2993
timestamp 1626908933
transform 1 0 11856 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1019
timestamp 1626908933
transform 1 0 12048 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2986
timestamp 1626908933
transform 1 0 12048 0 1 21645
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_116
timestamp 1626908933
transform 1 0 12480 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_473
timestamp 1626908933
transform 1 0 12480 0 -1 22644
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_199
timestamp 1626908933
transform 1 0 12500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_847
timestamp 1626908933
transform 1 0 12500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_199
timestamp 1626908933
transform 1 0 12500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_847
timestamp 1626908933
transform 1 0 12500 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_359
timestamp 1626908933
transform 1 0 12576 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_957
timestamp 1626908933
transform 1 0 12576 0 -1 22644
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3073
timestamp 1626908933
transform 1 0 12912 0 1 21497
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1138
timestamp 1626908933
transform 1 0 12912 0 1 21497
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3037
timestamp 1626908933
transform 1 0 13008 0 1 21497
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1070
timestamp 1626908933
transform 1 0 13008 0 1 21497
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3069
timestamp 1626908933
transform 1 0 12816 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1134
timestamp 1626908933
transform 1 0 12816 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3034
timestamp 1626908933
transform 1 0 12816 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1067
timestamp 1626908933
transform 1 0 12816 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3066
timestamp 1626908933
transform 1 0 13008 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1131
timestamp 1626908933
transform 1 0 13008 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3031
timestamp 1626908933
transform 1 0 13104 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1064
timestamp 1626908933
transform 1 0 13104 0 1 21645
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_458
timestamp 1626908933
transform 1 0 12960 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1180
timestamp 1626908933
transform 1 0 12960 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_723
timestamp 1626908933
transform 1 0 13728 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_122
timestamp 1626908933
transform 1 0 13728 0 -1 22644
box -38 -49 230 715
use L1M1_PR  L1M1_PR_3026
timestamp 1626908933
transform 1 0 13968 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1091
timestamp 1626908933
transform 1 0 13968 0 1 21423
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2992
timestamp 1626908933
transform 1 0 13872 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1025
timestamp 1626908933
transform 1 0 13872 0 1 21423
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1219
timestamp 1626908933
transform 1 0 13920 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_228
timestamp 1626908933
transform 1 0 13920 0 -1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3031
timestamp 1626908933
transform 1 0 14160 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1096
timestamp 1626908933
transform 1 0 14160 0 1 21867
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2998
timestamp 1626908933
transform 1 0 14160 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1031
timestamp 1626908933
transform 1 0 14160 0 1 21867
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2183
timestamp 1626908933
transform 1 0 14352 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_248
timestamp 1626908933
transform 1 0 14352 0 1 21867
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2195
timestamp 1626908933
transform 1 0 14352 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_228
timestamp 1626908933
transform 1 0 14352 0 1 21867
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_175
timestamp 1626908933
transform 1 0 14900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_823
timestamp 1626908933
transform 1 0 14900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_175
timestamp 1626908933
transform 1 0 14900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_823
timestamp 1626908933
transform 1 0 14900 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_427
timestamp 1626908933
transform 1 0 14016 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1149
timestamp 1626908933
transform 1 0 14016 0 -1 22644
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2201
timestamp 1626908933
transform 1 0 15216 0 1 22089
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2200
timestamp 1626908933
transform 1 0 16464 0 1 21793
box -29 -23 29 23
use L1M1_PR  L1M1_PR_266
timestamp 1626908933
transform 1 0 15216 0 1 22089
box -29 -23 29 23
use L1M1_PR  L1M1_PR_265
timestamp 1626908933
transform 1 0 16464 0 1 21793
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2211
timestamp 1626908933
transform 1 0 15216 0 1 21793
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2210
timestamp 1626908933
transform 1 0 15216 0 1 22089
box -32 -32 32 32
use M1M2_PR  M1M2_PR_244
timestamp 1626908933
transform 1 0 15216 0 1 21793
box -32 -32 32 32
use M1M2_PR  M1M2_PR_243
timestamp 1626908933
transform 1 0 15216 0 1 22089
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_79
timestamp 1626908933
transform -1 0 17472 0 -1 22644
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_33
timestamp 1626908933
transform -1 0 17472 0 -1 22644
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1050
timestamp 1626908933
transform 1 0 16656 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3017
timestamp 1626908933
transform 1 0 16656 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1117
timestamp 1626908933
transform 1 0 16848 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3052
timestamp 1626908933
transform 1 0 16848 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1116
timestamp 1626908933
transform 1 0 16656 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3051
timestamp 1626908933
transform 1 0 16656 0 1 21867
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1048
timestamp 1626908933
transform 1 0 16848 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3015
timestamp 1626908933
transform 1 0 16848 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1571
timestamp 1626908933
transform 1 0 17136 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3538
timestamp 1626908933
transform 1 0 17136 0 1 21867
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1660
timestamp 1626908933
transform 1 0 17040 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3595
timestamp 1626908933
transform 1 0 17040 0 1 21867
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_151
timestamp 1626908933
transform 1 0 17300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_799
timestamp 1626908933
transform 1 0 17300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_151
timestamp 1626908933
transform 1 0 17300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_799
timestamp 1626908933
transform 1 0 17300 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_115
timestamp 1626908933
transform 1 0 17472 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_472
timestamp 1626908933
transform 1 0 17472 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_227
timestamp 1626908933
transform 1 0 17568 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1218
timestamp 1626908933
transform 1 0 17568 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_226
timestamp 1626908933
transform 1 0 18048 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1217
timestamp 1626908933
transform 1 0 18048 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1535
timestamp 1626908933
transform 1 0 18192 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3502
timestamp 1626908933
transform 1 0 18192 0 1 21571
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_353
timestamp 1626908933
transform 1 0 18144 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1075
timestamp 1626908933
transform 1 0 18144 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_265
timestamp 1626908933
transform 1 0 17664 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_863
timestamp 1626908933
transform 1 0 17664 0 -1 22644
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1296
timestamp 1626908933
transform 1 0 18384 0 1 21497
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1394
timestamp 1626908933
transform 1 0 18480 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3231
timestamp 1626908933
transform 1 0 18384 0 1 21497
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3329
timestamp 1626908933
transform 1 0 18480 0 1 21645
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_121
timestamp 1626908933
transform 1 0 18912 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_722
timestamp 1626908933
transform 1 0 18912 0 -1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1309
timestamp 1626908933
transform 1 0 18864 0 1 21793
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3276
timestamp 1626908933
transform 1 0 18864 0 1 21793
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1295
timestamp 1626908933
transform 1 0 18768 0 1 21497
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1390
timestamp 1626908933
transform 1 0 18960 0 1 21793
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3230
timestamp 1626908933
transform 1 0 18768 0 1 21497
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3325
timestamp 1626908933
transform 1 0 18960 0 1 21793
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_238
timestamp 1626908933
transform 1 0 19104 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_836
timestamp 1626908933
transform 1 0 19104 0 -1 22644
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1432
timestamp 1626908933
transform 1 0 19632 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3399
timestamp 1626908933
transform 1 0 19632 0 1 21571
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1518
timestamp 1626908933
transform 1 0 19632 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3453
timestamp 1626908933
transform 1 0 19632 0 1 21571
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1312
timestamp 1626908933
transform 1 0 20112 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3279
timestamp 1626908933
transform 1 0 20112 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1394
timestamp 1626908933
transform 1 0 20304 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3361
timestamp 1626908933
transform 1 0 20304 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1478
timestamp 1626908933
transform 1 0 20304 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3413
timestamp 1626908933
transform 1 0 20304 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1532
timestamp 1626908933
transform 1 0 20400 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3499
timestamp 1626908933
transform 1 0 20400 0 1 21571
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1620
timestamp 1626908933
transform 1 0 21264 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3555
timestamp 1626908933
transform 1 0 21264 0 1 21571
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_127
timestamp 1626908933
transform 1 0 19700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_775
timestamp 1626908933
transform 1 0 19700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_127
timestamp 1626908933
transform 1 0 19700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_775
timestamp 1626908933
transform 1 0 19700 0 1 21978
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1385
timestamp 1626908933
transform 1 0 21648 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3352
timestamp 1626908933
transform 1 0 21648 0 1 21867
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1467
timestamp 1626908933
transform 1 0 21648 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3402
timestamp 1626908933
transform 1 0 21648 0 1 21867
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_103
timestamp 1626908933
transform 1 0 22100 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_751
timestamp 1626908933
transform 1 0 22100 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_103
timestamp 1626908933
transform 1 0 22100 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_751
timestamp 1626908933
transform 1 0 22100 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_59
timestamp 1626908933
transform -1 0 22176 0 -1 22644
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_13
timestamp 1626908933
transform -1 0 22176 0 -1 22644
box -38 -49 2726 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_114
timestamp 1626908933
transform 1 0 22464 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_471
timestamp 1626908933
transform 1 0 22464 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_543
timestamp 1626908933
transform 1 0 22176 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1144
timestamp 1626908933
transform 1 0 22176 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_913
timestamp 1626908933
transform 1 0 22368 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1904
timestamp 1626908933
transform 1 0 22368 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1838
timestamp 1626908933
transform 1 0 22320 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3805
timestamp 1626908933
transform 1 0 22320 0 1 21645
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_914
timestamp 1626908933
transform 1 0 22560 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1905
timestamp 1626908933
transform 1 0 22560 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_4
timestamp 1626908933
transform -1 0 23424 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_10
timestamp 1626908933
transform -1 0 23424 0 -1 22644
box -38 -49 806 715
use L1M1_PR  L1M1_PR_393
timestamp 1626908933
transform 1 0 23184 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1820
timestamp 1626908933
transform 1 0 23184 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2328
timestamp 1626908933
transform 1 0 23184 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3755
timestamp 1626908933
transform 1 0 23184 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3803
timestamp 1626908933
transform 1 0 23568 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2350
timestamp 1626908933
transform 1 0 23472 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1868
timestamp 1626908933
transform 1 0 23568 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_415
timestamp 1626908933
transform 1 0 23472 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3736
timestamp 1626908933
transform 1 0 23760 0 1 21571
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1801
timestamp 1626908933
transform 1 0 23760 0 1 21571
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1906
timestamp 1626908933
transform 1 0 23616 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_915
timestamp 1626908933
transform 1 0 23616 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1145
timestamp 1626908933
transform 1 0 23424 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_544
timestamp 1626908933
transform 1 0 23424 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_5
timestamp 1626908933
transform -1 0 24480 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_11
timestamp 1626908933
transform -1 0 24480 0 -1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_369
timestamp 1626908933
transform 1 0 24144 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1898
timestamp 1626908933
transform 1 0 24048 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2336
timestamp 1626908933
transform 1 0 24144 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3865
timestamp 1626908933
transform 1 0 24048 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_419
timestamp 1626908933
transform 1 0 24240 0 1 21793
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2386
timestamp 1626908933
transform 1 0 24240 0 1 21793
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_79
timestamp 1626908933
transform 1 0 24500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_727
timestamp 1626908933
transform 1 0 24500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_79
timestamp 1626908933
transform 1 0 24500 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_727
timestamp 1626908933
transform 1 0 24500 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_200
timestamp 1626908933
transform 1 0 24480 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_922
timestamp 1626908933
transform 1 0 24480 0 -1 22644
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1492
timestamp 1626908933
transform 1 0 25104 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3427
timestamp 1626908933
transform 1 0 25104 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1378
timestamp 1626908933
transform 1 0 25488 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1409
timestamp 1626908933
transform 1 0 25392 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3345
timestamp 1626908933
transform 1 0 25488 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3376
timestamp 1626908933
transform 1 0 25392 0 1 21645
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1458
timestamp 1626908933
transform 1 0 25488 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3393
timestamp 1626908933
transform 1 0 25488 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1803
timestamp 1626908933
transform 1 0 26256 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3770
timestamp 1626908933
transform 1 0 26256 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_381
timestamp 1626908933
transform 1 0 26544 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2348
timestamp 1626908933
transform 1 0 26544 0 1 21645
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_83
timestamp 1626908933
transform 1 0 27072 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_681
timestamp 1626908933
transform 1 0 27072 0 -1 22644
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_55
timestamp 1626908933
transform 1 0 26900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_703
timestamp 1626908933
transform 1 0 26900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_55
timestamp 1626908933
transform 1 0 26900 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_703
timestamp 1626908933
transform 1 0 26900 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_113
timestamp 1626908933
transform 1 0 27456 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_470
timestamp 1626908933
transform 1 0 27456 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_120
timestamp 1626908933
transform 1 0 27552 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_721
timestamp 1626908933
transform 1 0 27552 0 -1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_352
timestamp 1626908933
transform 1 0 27312 0 1 21867
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2319
timestamp 1626908933
transform 1 0 27312 0 1 21867
box -32 -32 32 32
use L1M1_PR  L1M1_PR_374
timestamp 1626908933
transform 1 0 27312 0 1 21867
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2309
timestamp 1626908933
transform 1 0 27312 0 1 21867
box -29 -23 29 23
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_18
timestamp 1626908933
transform -1 0 27072 0 -1 22644
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_6
timestamp 1626908933
transform -1 0 27072 0 -1 22644
box -38 -49 1862 715
use M1M2_PR  M1M2_PR_2384
timestamp 1626908933
transform 1 0 27888 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_417
timestamp 1626908933
transform 1 0 27888 0 1 21571
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_843
timestamp 1626908933
transform 1 0 27744 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_121
timestamp 1626908933
transform 1 0 27744 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_916
timestamp 1626908933
transform 1 0 28512 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1907
timestamp 1626908933
transform 1 0 28512 0 -1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_373
timestamp 1626908933
transform 1 0 28560 0 1 21793
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1814
timestamp 1626908933
transform 1 0 28752 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2308
timestamp 1626908933
transform 1 0 28560 0 1 21793
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3749
timestamp 1626908933
transform 1 0 28752 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3730
timestamp 1626908933
transform 1 0 29232 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1795
timestamp 1626908933
transform 1 0 29232 0 1 21423
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3798
timestamp 1626908933
transform 1 0 29040 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2345
timestamp 1626908933
transform 1 0 28944 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1863
timestamp 1626908933
transform 1 0 29040 0 1 21645
box -29 -23 29 23
use L1M1_PR  L1M1_PR_410
timestamp 1626908933
transform 1 0 28944 0 1 21645
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3857
timestamp 1626908933
transform 1 0 29040 0 1 21645
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1890
timestamp 1626908933
transform 1 0 29040 0 1 21645
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_679
timestamp 1626908933
transform 1 0 29300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_31
timestamp 1626908933
transform 1 0 29300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_679
timestamp 1626908933
transform 1 0 29300 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_31
timestamp 1626908933
transform 1 0 29300 0 1 21978
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3729
timestamp 1626908933
transform 1 0 29232 0 1 22089
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1794
timestamp 1626908933
transform 1 0 29232 0 1 22089
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3751
timestamp 1626908933
transform 1 0 29136 0 1 22089
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1784
timestamp 1626908933
transform 1 0 29136 0 1 22089
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_40
timestamp 1626908933
transform 1 0 29280 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_638
timestamp 1626908933
transform 1 0 29280 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_8
timestamp 1626908933
transform 1 0 28608 0 -1 22644
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_23
timestamp 1626908933
transform 1 0 28608 0 -1 22644
box -38 -49 710 715
use M1M2_PR  M1M2_PR_3754
timestamp 1626908933
transform 1 0 29616 0 1 21423
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1787
timestamp 1626908933
transform 1 0 29616 0 1 21423
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_794
timestamp 1626908933
transform 1 0 29664 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_72
timestamp 1626908933
transform 1 0 29664 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_225
timestamp 1626908933
transform 1 0 30432 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1216
timestamp 1626908933
transform 1 0 30432 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_409
timestamp 1626908933
transform 1 0 30672 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2376
timestamp 1626908933
transform 1 0 30672 0 1 21571
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1823
timestamp 1626908933
transform 1 0 31248 0 1 21719
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3790
timestamp 1626908933
transform 1 0 31248 0 1 21719
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_26
timestamp 1626908933
transform 1 0 30912 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_748
timestamp 1626908933
transform 1 0 30912 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_20
timestamp 1626908933
transform 1 0 30528 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_618
timestamp 1626908933
transform 1 0 30528 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_112
timestamp 1626908933
transform 1 0 31680 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_469
timestamp 1626908933
transform 1 0 31680 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_545
timestamp 1626908933
transform 1 0 31776 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1146
timestamp 1626908933
transform 1 0 31776 0 -1 22644
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_7
timestamp 1626908933
transform 1 0 31700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_655
timestamp 1626908933
transform 1 0 31700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_7
timestamp 1626908933
transform 1 0 31700 0 1 21978
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_655
timestamp 1626908933
transform 1 0 31700 0 1 21978
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_917
timestamp 1626908933
transform 1 0 31968 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1908
timestamp 1626908933
transform 1 0 31968 0 -1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3815
timestamp 1626908933
transform 1 0 48 0 1 22903
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1848
timestamp 1626908933
transform 1 0 48 0 1 22903
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1909
timestamp 1626908933
transform 1 0 192 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_918
timestamp 1626908933
transform 1 0 192 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_468
timestamp 1626908933
transform 1 0 288 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_111
timestamp 1626908933
transform 1 0 288 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1147
timestamp 1626908933
transform 1 0 0 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_546
timestamp 1626908933
transform 1 0 0 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1189
timestamp 1626908933
transform 1 0 384 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_591
timestamp 1626908933
transform 1 0 384 0 1 22644
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1279
timestamp 1626908933
transform 1 0 1700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_631
timestamp 1626908933
transform 1 0 1700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1279
timestamp 1626908933
transform 1 0 1700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_631
timestamp 1626908933
transform 1 0 1700 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_61
timestamp 1626908933
transform -1 0 3456 0 1 22644
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_15
timestamp 1626908933
transform -1 0 3456 0 1 22644
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3118
timestamp 1626908933
transform 1 0 3408 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1183
timestamp 1626908933
transform 1 0 3408 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3081
timestamp 1626908933
transform 1 0 3312 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1114
timestamp 1626908933
transform 1 0 3312 0 1 22311
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2247
timestamp 1626908933
transform 1 0 3024 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_312
timestamp 1626908933
transform 1 0 3024 0 1 22533
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2258
timestamp 1626908933
transform 1 0 2928 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_291
timestamp 1626908933
transform 1 0 2928 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3514
timestamp 1626908933
transform 1 0 3408 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1547
timestamp 1626908933
transform 1 0 3408 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3570
timestamp 1626908933
transform 1 0 3600 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1635
timestamp 1626908933
transform 1 0 3600 0 1 22533
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_626
timestamp 1626908933
transform 1 0 3456 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1348
timestamp 1626908933
transform 1 0 3456 0 1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_471
timestamp 1626908933
transform 1 0 4272 0 1 22829
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2438
timestamp 1626908933
transform 1 0 4272 0 1 22829
box -32 -32 32 32
use L1M1_PR  L1M1_PR_469
timestamp 1626908933
transform 1 0 4176 0 1 22829
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2404
timestamp 1626908933
transform 1 0 4176 0 1 22829
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_607
timestamp 1626908933
transform 1 0 4100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1255
timestamp 1626908933
transform 1 0 4100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_607
timestamp 1626908933
transform 1 0 4100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1255
timestamp 1626908933
transform 1 0 4100 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_55
timestamp 1626908933
transform 1 0 4224 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_117
timestamp 1626908933
transform 1 0 4224 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1910
timestamp 1626908933
transform 1 0 5280 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_919
timestamp 1626908933
transform 1 0 5280 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1148
timestamp 1626908933
transform 1 0 5088 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_547
timestamp 1626908933
transform 1 0 5088 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_98
timestamp 1626908933
transform 1 0 4608 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_46
timestamp 1626908933
transform 1 0 4608 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_467
timestamp 1626908933
transform 1 0 4992 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_110
timestamp 1626908933
transform 1 0 4992 0 1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2444
timestamp 1626908933
transform 1 0 5520 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_509
timestamp 1626908933
transform 1 0 5520 0 1 22755
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2481
timestamp 1626908933
transform 1 0 5424 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2480
timestamp 1626908933
transform 1 0 5424 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_514
timestamp 1626908933
transform 1 0 5424 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_513
timestamp 1626908933
transform 1 0 5424 0 1 22755
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_58
timestamp 1626908933
transform -1 0 5856 0 1 22644
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_127
timestamp 1626908933
transform -1 0 5856 0 1 22644
box -38 -49 518 715
use L1M1_PR  L1M1_PR_2443
timestamp 1626908933
transform 1 0 5616 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_508
timestamp 1626908933
transform 1 0 5616 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3179
timestamp 1626908933
transform 1 0 5712 0 1 22163
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2450
timestamp 1626908933
transform 1 0 5808 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1244
timestamp 1626908933
transform 1 0 5712 0 1 22163
box -29 -23 29 23
use L1M1_PR  L1M1_PR_515
timestamp 1626908933
transform 1 0 5808 0 1 22385
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2486
timestamp 1626908933
transform 1 0 5808 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_519
timestamp 1626908933
transform 1 0 5808 0 1 22385
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1215
timestamp 1626908933
transform 1 0 5856 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_224
timestamp 1626908933
transform 1 0 5856 0 1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3181
timestamp 1626908933
transform 1 0 5904 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1246
timestamp 1626908933
transform 1 0 5904 0 1 22385
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3151
timestamp 1626908933
transform 1 0 6096 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1184
timestamp 1626908933
transform 1 0 6096 0 1 22385
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3768
timestamp 1626908933
transform 1 0 6000 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1833
timestamp 1626908933
transform 1 0 6000 0 1 22533
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3824
timestamp 1626908933
transform 1 0 6000 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1857
timestamp 1626908933
transform 1 0 6000 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2447
timestamp 1626908933
transform 1 0 6288 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_512
timestamp 1626908933
transform 1 0 6288 0 1 22533
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2484
timestamp 1626908933
transform 1 0 6288 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_517
timestamp 1626908933
transform 1 0 6288 0 1 22533
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_590
timestamp 1626908933
transform 1 0 5952 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1312
timestamp 1626908933
transform 1 0 5952 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_223
timestamp 1626908933
transform 1 0 6720 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1214
timestamp 1626908933
transform 1 0 6720 0 1 22644
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_583
timestamp 1626908933
transform 1 0 6500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1231
timestamp 1626908933
transform 1 0 6500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_583
timestamp 1626908933
transform 1 0 6500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1231
timestamp 1626908933
transform 1 0 6500 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_566
timestamp 1626908933
transform 1 0 7200 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1288
timestamp 1626908933
transform 1 0 7200 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_479
timestamp 1626908933
transform 1 0 6816 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1077
timestamp 1626908933
transform 1 0 6816 0 1 22644
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3196
timestamp 1626908933
transform 1 0 7824 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2230
timestamp 1626908933
transform 1 0 7920 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1261
timestamp 1626908933
transform 1 0 7824 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_295
timestamp 1626908933
transform 1 0 7920 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2241
timestamp 1626908933
transform 1 0 7920 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_274
timestamp 1626908933
transform 1 0 7920 0 1 22311
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3180
timestamp 1626908933
transform 1 0 7632 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1245
timestamp 1626908933
transform 1 0 7632 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3186
timestamp 1626908933
transform 1 0 7920 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1251
timestamp 1626908933
transform 1 0 7920 0 1 22533
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_458
timestamp 1626908933
transform 1 0 7968 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1056
timestamp 1626908933
transform 1 0 7968 0 1 22644
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2416
timestamp 1626908933
transform 1 0 8208 0 1 22237
box -29 -23 29 23
use L1M1_PR  L1M1_PR_481
timestamp 1626908933
transform 1 0 8208 0 1 22237
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3165
timestamp 1626908933
transform 1 0 8112 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1198
timestamp 1626908933
transform 1 0 8112 0 1 22237
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_222
timestamp 1626908933
transform 1 0 8352 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1213
timestamp 1626908933
transform 1 0 8352 0 1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1189
timestamp 1626908933
transform 1 0 8688 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3156
timestamp 1626908933
transform 1 0 8688 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_294
timestamp 1626908933
transform 1 0 8880 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1164
timestamp 1626908933
transform 1 0 9072 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2229
timestamp 1626908933
transform 1 0 8880 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3099
timestamp 1626908933
transform 1 0 9072 0 1 22533
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_559
timestamp 1626908933
transform 1 0 8900 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1207
timestamp 1626908933
transform 1 0 8900 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_559
timestamp 1626908933
transform 1 0 8900 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1207
timestamp 1626908933
transform 1 0 8900 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_547
timestamp 1626908933
transform 1 0 8448 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1269
timestamp 1626908933
transform 1 0 8448 0 1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1096
timestamp 1626908933
transform 1 0 9264 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3063
timestamp 1626908933
transform 1 0 9264 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1160
timestamp 1626908933
transform 1 0 9264 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3095
timestamp 1626908933
transform 1 0 9264 0 1 22385
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_109
timestamp 1626908933
transform 1 0 9984 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_466
timestamp 1626908933
transform 1 0 9984 0 1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_480
timestamp 1626908933
transform 1 0 9840 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1092
timestamp 1626908933
transform 1 0 9840 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2447
timestamp 1626908933
transform 1 0 9840 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3059
timestamp 1626908933
transform 1 0 9840 0 1 22385
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_524
timestamp 1626908933
transform 1 0 9216 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1246
timestamp 1626908933
transform 1 0 9216 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1017
timestamp 1626908933
transform 1 0 10080 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_419
timestamp 1626908933
transform 1 0 10080 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1232
timestamp 1626908933
transform 1 0 10464 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_510
timestamp 1626908933
transform 1 0 10464 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_221
timestamp 1626908933
transform 1 0 11232 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1212
timestamp 1626908933
transform 1 0 11232 0 1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_479
timestamp 1626908933
transform 1 0 11472 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2446
timestamp 1626908933
transform 1 0 11472 0 1 22311
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_535
timestamp 1626908933
transform 1 0 11300 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1183
timestamp 1626908933
transform 1 0 11300 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_535
timestamp 1626908933
transform 1 0 11300 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1183
timestamp 1626908933
transform 1 0 11300 0 1 22644
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1587
timestamp 1626908933
transform 1 0 11856 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3554
timestamp 1626908933
transform 1 0 11856 0 1 22385
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_479
timestamp 1626908933
transform 1 0 11712 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1201
timestamp 1626908933
transform 1 0 11712 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_392
timestamp 1626908933
transform 1 0 11328 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_990
timestamp 1626908933
transform 1 0 11328 0 1 22644
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3645
timestamp 1626908933
transform 1 0 12048 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3610
timestamp 1626908933
transform 1 0 12432 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1710
timestamp 1626908933
transform 1 0 12048 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1675
timestamp 1626908933
transform 1 0 12432 0 1 22385
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3585
timestamp 1626908933
transform 1 0 12624 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1618
timestamp 1626908933
transform 1 0 12624 0 1 22311
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_968
timestamp 1626908933
transform 1 0 12480 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_370
timestamp 1626908933
transform 1 0 12480 0 1 22644
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3689
timestamp 1626908933
transform 1 0 13488 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1722
timestamp 1626908933
transform 1 0 13488 0 1 22237
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1211
timestamp 1626908933
transform 1 0 12864 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_220
timestamp 1626908933
transform 1 0 12864 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1179
timestamp 1626908933
transform 1 0 12960 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_457
timestamp 1626908933
transform 1 0 12960 0 1 22644
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1159
timestamp 1626908933
transform 1 0 13700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_511
timestamp 1626908933
transform 1 0 13700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1159
timestamp 1626908933
transform 1 0 13700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_511
timestamp 1626908933
transform 1 0 13700 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_67
timestamp 1626908933
transform -1 0 14304 0 1 22644
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_28
timestamp 1626908933
transform -1 0 14304 0 1 22644
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2185
timestamp 1626908933
transform 1 0 13680 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_250
timestamp 1626908933
transform 1 0 13680 0 1 22755
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_341
timestamp 1626908933
transform 1 0 14304 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_939
timestamp 1626908933
transform 1 0 14304 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_548
timestamp 1626908933
transform 1 0 14688 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1149
timestamp 1626908933
transform 1 0 14688 0 1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_227
timestamp 1626908933
transform 1 0 14352 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1609
timestamp 1626908933
transform 1 0 14640 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2194
timestamp 1626908933
transform 1 0 14352 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3576
timestamp 1626908933
transform 1 0 14640 0 1 22385
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_108
timestamp 1626908933
transform 1 0 14976 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_465
timestamp 1626908933
transform 1 0 14976 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_549
timestamp 1626908933
transform 1 0 15072 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1150
timestamp 1626908933
transform 1 0 15072 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_920
timestamp 1626908933
transform 1 0 14880 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1911
timestamp 1626908933
transform 1 0 14880 0 1 22644
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1135
timestamp 1626908933
transform 1 0 16100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_487
timestamp 1626908933
transform 1 0 16100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1135
timestamp 1626908933
transform 1 0 16100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_487
timestamp 1626908933
transform 1 0 16100 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_90
timestamp 1626908933
transform -1 0 17952 0 1 22644
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_44
timestamp 1626908933
transform -1 0 17952 0 1 22644
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3635
timestamp 1626908933
transform 1 0 17040 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3594
timestamp 1626908933
transform 1 0 17424 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1700
timestamp 1626908933
transform 1 0 17040 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1659
timestamp 1626908933
transform 1 0 17424 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3676
timestamp 1626908933
transform 1 0 16656 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3537
timestamp 1626908933
transform 1 0 17136 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1709
timestamp 1626908933
transform 1 0 16656 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1570
timestamp 1626908933
transform 1 0 17136 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3571
timestamp 1626908933
transform 1 0 17520 0 1 22459
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1604
timestamp 1626908933
transform 1 0 17520 0 1 22459
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1210
timestamp 1626908933
transform 1 0 17952 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_219
timestamp 1626908933
transform 1 0 17952 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1074
timestamp 1626908933
transform 1 0 18048 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_352
timestamp 1626908933
transform 1 0 18048 0 1 22644
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1111
timestamp 1626908933
transform 1 0 18500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_463
timestamp 1626908933
transform 1 0 18500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1111
timestamp 1626908933
transform 1 0 18500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_463
timestamp 1626908933
transform 1 0 18500 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_9
timestamp 1626908933
transform 1 0 18816 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_3
timestamp 1626908933
transform 1 0 18816 0 1 22644
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3760
timestamp 1626908933
transform 1 0 18864 0 1 22903
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1825
timestamp 1626908933
transform 1 0 18864 0 1 22903
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2361
timestamp 1626908933
transform 1 0 19152 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_394
timestamp 1626908933
transform 1 0 19152 0 1 22237
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_107
timestamp 1626908933
transform 1 0 19968 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_464
timestamp 1626908933
transform 1 0 19968 0 1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_336
timestamp 1626908933
transform 1 0 19920 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2303
timestamp 1626908933
transform 1 0 19920 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_360
timestamp 1626908933
transform 1 0 19824 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2295
timestamp 1626908933
transform 1 0 19824 0 1 22533
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_306
timestamp 1626908933
transform 1 0 20064 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1028
timestamp 1626908933
transform 1 0 20064 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_220
timestamp 1626908933
transform 1 0 19584 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_818
timestamp 1626908933
transform 1 0 19584 0 1 22644
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1361
timestamp 1626908933
transform 1 0 20208 0 1 22903
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3328
timestamp 1626908933
transform 1 0 20208 0 1 22903
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1443
timestamp 1626908933
transform 1 0 20880 0 1 22903
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3378
timestamp 1626908933
transform 1 0 20880 0 1 22903
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_439
timestamp 1626908933
transform 1 0 20900 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1087
timestamp 1626908933
transform 1 0 20900 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_439
timestamp 1626908933
transform 1 0 20900 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1087
timestamp 1626908933
transform 1 0 20900 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_17
timestamp 1626908933
transform 1 0 20832 0 1 22644
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_42
timestamp 1626908933
transform 1 0 20832 0 1 22644
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1384
timestamp 1626908933
transform 1 0 21648 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1417
timestamp 1626908933
transform 1 0 21264 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3351
timestamp 1626908933
transform 1 0 21648 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3384
timestamp 1626908933
transform 1 0 21264 0 1 22385
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1466
timestamp 1626908933
transform 1 0 21744 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3401
timestamp 1626908933
transform 1 0 21744 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1416
timestamp 1626908933
transform 1 0 21264 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1428
timestamp 1626908933
transform 1 0 21456 0 1 22903
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3383
timestamp 1626908933
transform 1 0 21264 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3395
timestamp 1626908933
transform 1 0 21456 0 1 22903
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1502
timestamp 1626908933
transform 1 0 21168 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1515
timestamp 1626908933
transform 1 0 21072 0 1 22903
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3437
timestamp 1626908933
transform 1 0 21168 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3450
timestamp 1626908933
transform 1 0 21072 0 1 22903
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_281
timestamp 1626908933
transform 1 0 21312 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1003
timestamp 1626908933
transform 1 0 21312 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_782
timestamp 1626908933
transform 1 0 22080 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_184
timestamp 1626908933
transform 1 0 22080 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_921
timestamp 1626908933
transform 1 0 22464 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1912
timestamp 1626908933
transform 1 0 22464 0 1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1501
timestamp 1626908933
transform 1 0 22128 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3436
timestamp 1626908933
transform 1 0 22128 0 1 22385
box -29 -23 29 23
use M1M2_PR  M1M2_PR_333
timestamp 1626908933
transform 1 0 22608 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2300
timestamp 1626908933
transform 1 0 22608 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1233
timestamp 1626908933
transform 1 0 22896 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3168
timestamp 1626908933
transform 1 0 22896 0 1 22533
box -29 -23 29 23
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_1
timestamp 1626908933
transform -1 0 23040 0 1 22644
box -38 -49 518 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_3
timestamp 1626908933
transform -1 0 23040 0 1 22644
box -38 -49 518 715
use L1M1_PR  L1M1_PR_3292
timestamp 1626908933
transform 1 0 23088 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1357
timestamp 1626908933
transform 1 0 23088 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3236
timestamp 1626908933
transform 1 0 23088 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3129
timestamp 1626908933
transform 1 0 22992 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1269
timestamp 1626908933
transform 1 0 23088 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1162
timestamp 1626908933
transform 1 0 22992 0 1 22533
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1063
timestamp 1626908933
transform 1 0 23300 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_415
timestamp 1626908933
transform 1 0 23300 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1063
timestamp 1626908933
transform 1 0 23300 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_415
timestamp 1626908933
transform 1 0 23300 0 1 22644
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3167
timestamp 1626908933
transform 1 0 22992 0 1 22903
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1232
timestamp 1626908933
transform 1 0 22992 0 1 22903
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3128
timestamp 1626908933
transform 1 0 22992 0 1 22903
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1161
timestamp 1626908933
transform 1 0 22992 0 1 22903
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_720
timestamp 1626908933
transform 1 0 23040 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_119
timestamp 1626908933
transform 1 0 23040 0 1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1302
timestamp 1626908933
transform 1 0 23472 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3269
timestamp 1626908933
transform 1 0 23472 0 1 22311
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_231
timestamp 1626908933
transform 1 0 23232 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_953
timestamp 1626908933
transform 1 0 23232 0 1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_373
timestamp 1626908933
transform 1 0 24336 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1897
timestamp 1626908933
transform 1 0 24048 0 1 22459
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2340
timestamp 1626908933
transform 1 0 24336 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3864
timestamp 1626908933
transform 1 0 24048 0 1 22459
box -32 -32 32 32
use L1M1_PR  L1M1_PR_395
timestamp 1626908933
transform 1 0 24432 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1385
timestamp 1626908933
transform 1 0 23952 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2330
timestamp 1626908933
transform 1 0 24432 0 1 22385
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3320
timestamp 1626908933
transform 1 0 23952 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_372
timestamp 1626908933
transform 1 0 24336 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1896
timestamp 1626908933
transform 1 0 24048 0 1 22903
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2339
timestamp 1626908933
transform 1 0 24336 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3863
timestamp 1626908933
transform 1 0 24048 0 1 22903
box -32 -32 32 32
use L1M1_PR  L1M1_PR_396
timestamp 1626908933
transform 1 0 24048 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2331
timestamp 1626908933
transform 1 0 24048 0 1 22755
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_0
timestamp 1626908933
transform 1 0 24000 0 1 22644
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_15
timestamp 1626908933
transform 1 0 24000 0 1 22644
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1913
timestamp 1626908933
transform 1 0 24864 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_922
timestamp 1626908933
transform 1 0 24864 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1151
timestamp 1626908933
transform 1 0 24672 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_550
timestamp 1626908933
transform 1 0 24672 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_106
timestamp 1626908933
transform 1 0 24960 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_463
timestamp 1626908933
transform 1 0 24960 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_218
timestamp 1626908933
transform 1 0 25056 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1209
timestamp 1626908933
transform 1 0 25056 0 1 22644
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1434
timestamp 1626908933
transform 1 0 25392 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3369
timestamp 1626908933
transform 1 0 25392 0 1 22533
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_391
timestamp 1626908933
transform 1 0 25700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1039
timestamp 1626908933
transform 1 0 25700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_391
timestamp 1626908933
transform 1 0 25700 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1039
timestamp 1626908933
transform 1 0 25700 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_181
timestamp 1626908933
transform 1 0 25152 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_903
timestamp 1626908933
transform 1 0 25152 0 1 22644
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3304
timestamp 1626908933
transform 1 0 25776 0 1 22237
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1369
timestamp 1626908933
transform 1 0 25776 0 1 22237
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3244
timestamp 1626908933
transform 1 0 26064 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1277
timestamp 1626908933
transform 1 0 26064 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3318
timestamp 1626908933
transform 1 0 25872 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1351
timestamp 1626908933
transform 1 0 25872 0 1 22533
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3368
timestamp 1626908933
transform 1 0 25872 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1433
timestamp 1626908933
transform 1 0 25872 0 1 22755
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3317
timestamp 1626908933
transform 1 0 25872 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1350
timestamp 1626908933
transform 1 0 25872 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3388
timestamp 1626908933
transform 1 0 26064 0 1 22903
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1421
timestamp 1626908933
transform 1 0 26064 0 1 22903
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3442
timestamp 1626908933
transform 1 0 26160 0 1 22903
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1507
timestamp 1626908933
transform 1 0 26160 0 1 22903
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3305
timestamp 1626908933
transform 1 0 26352 0 1 22237
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1370
timestamp 1626908933
transform 1 0 26352 0 1 22237
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3247
timestamp 1626908933
transform 1 0 26352 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1280
timestamp 1626908933
transform 1 0 26352 0 1 22237
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1208
timestamp 1626908933
transform 1 0 26400 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_217
timestamp 1626908933
transform 1 0 26400 0 1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2305
timestamp 1626908933
transform 1 0 26544 0 1 22755
box -32 -32 32 32
use M1M2_PR  M1M2_PR_338
timestamp 1626908933
transform 1 0 26544 0 1 22755
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_152
timestamp 1626908933
transform 1 0 26496 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_874
timestamp 1626908933
transform 1 0 26496 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_15
timestamp 1626908933
transform 1 0 25920 0 1 22644
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_40
timestamp 1626908933
transform 1 0 25920 0 1 22644
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1299
timestamp 1626908933
transform 1 0 26736 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3266
timestamp 1626908933
transform 1 0 26736 0 1 22311
box -32 -32 32 32
use L1M1_PR  L1M1_PR_375
timestamp 1626908933
transform 1 0 26928 0 1 22237
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2310
timestamp 1626908933
transform 1 0 26928 0 1 22237
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_216
timestamp 1626908933
transform 1 0 27264 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1207
timestamp 1626908933
transform 1 0 27264 0 1 22644
box -38 -49 134 715
use M1M2_PR  M1M2_PR_348
timestamp 1626908933
transform 1 0 27408 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_351
timestamp 1626908933
transform 1 0 27312 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2315
timestamp 1626908933
transform 1 0 27408 0 1 22533
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2318
timestamp 1626908933
transform 1 0 27312 0 1 22237
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_82
timestamp 1626908933
transform 1 0 27360 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_680
timestamp 1626908933
transform 1 0 27360 0 1 22644
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2383
timestamp 1626908933
transform 1 0 27888 0 1 22237
box -32 -32 32 32
use M1M2_PR  M1M2_PR_416
timestamp 1626908933
transform 1 0 27888 0 1 22237
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1015
timestamp 1626908933
transform 1 0 28100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_367
timestamp 1626908933
transform 1 0 28100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1015
timestamp 1626908933
transform 1 0 28100 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_367
timestamp 1626908933
transform 1 0 28100 0 1 22644
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3745
timestamp 1626908933
transform 1 0 27888 0 1 22829
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2296
timestamp 1626908933
transform 1 0 27984 0 1 22755
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1810
timestamp 1626908933
transform 1 0 27888 0 1 22829
box -29 -23 29 23
use L1M1_PR  L1M1_PR_361
timestamp 1626908933
transform 1 0 27984 0 1 22755
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_719
timestamp 1626908933
transform 1 0 27744 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_118
timestamp 1626908933
transform 1 0 27744 0 1 22644
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1893
timestamp 1626908933
transform 1 0 28368 0 1 22385
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3860
timestamp 1626908933
transform 1 0 28368 0 1 22385
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_11
timestamp 1626908933
transform 1 0 27936 0 1 22644
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_26
timestamp 1626908933
transform 1 0 27936 0 1 22644
box -38 -49 710 715
use M1M2_PR  M1M2_PR_3787
timestamp 1626908933
transform 1 0 28560 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1820
timestamp 1626908933
transform 1 0 28560 0 1 22311
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3748
timestamp 1626908933
transform 1 0 28656 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1813
timestamp 1626908933
transform 1 0 28656 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2344
timestamp 1626908933
transform 1 0 28944 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_409
timestamp 1626908933
transform 1 0 28944 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3797
timestamp 1626908933
transform 1 0 29040 0 1 22311
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1862
timestamp 1626908933
transform 1 0 29040 0 1 22311
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3856
timestamp 1626908933
transform 1 0 29040 0 1 22311
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1889
timestamp 1626908933
transform 1 0 29040 0 1 22311
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2305
timestamp 1626908933
transform 1 0 28656 0 1 22533
box -29 -23 29 23
use L1M1_PR  L1M1_PR_370
timestamp 1626908933
transform 1 0 28656 0 1 22533
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_87
timestamp 1626908933
transform 1 0 28992 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_809
timestamp 1626908933
transform 1 0 28992 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_48
timestamp 1626908933
transform 1 0 28608 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_646
timestamp 1626908933
transform 1 0 28608 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1152
timestamp 1626908933
transform 1 0 29760 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_718
timestamp 1626908933
transform 1 0 30048 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_551
timestamp 1626908933
transform 1 0 29760 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_117
timestamp 1626908933
transform 1 0 30048 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_462
timestamp 1626908933
transform 1 0 29952 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_105
timestamp 1626908933
transform 1 0 29952 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1206
timestamp 1626908933
transform 1 0 30240 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_215
timestamp 1626908933
transform 1 0 30240 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_762
timestamp 1626908933
transform 1 0 30336 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_40
timestamp 1626908933
transform 1 0 30336 0 1 22644
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_991
timestamp 1626908933
transform 1 0 30500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_343
timestamp 1626908933
transform 1 0 30500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_991
timestamp 1626908933
transform 1 0 30500 0 1 22644
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_343
timestamp 1626908933
transform 1 0 30500 0 1 22644
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1205
timestamp 1626908933
transform 1 0 31104 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_214
timestamp 1626908933
transform 1 0 31104 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_728
timestamp 1626908933
transform 1 0 31200 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_6
timestamp 1626908933
transform 1 0 31200 0 1 22644
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3782
timestamp 1626908933
transform 1 0 31632 0 1 22829
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1815
timestamp 1626908933
transform 1 0 31632 0 1 22829
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1914
timestamp 1626908933
transform 1 0 31968 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_923
timestamp 1626908933
transform 1 0 31968 0 1 22644
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_966
timestamp 1626908933
transform 1 0 500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_318
timestamp 1626908933
transform 1 0 500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_966
timestamp 1626908933
transform 1 0 500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_318
timestamp 1626908933
transform 1 0 500 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_717
timestamp 1626908933
transform 1 0 0 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_116
timestamp 1626908933
transform 1 0 0 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1428
timestamp 1626908933
transform 1 0 192 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_706
timestamp 1626908933
transform 1 0 192 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_213
timestamp 1626908933
transform 1 0 960 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1204
timestamp 1626908933
transform 1 0 960 0 -1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_313
timestamp 1626908933
transform 1 0 1200 0 1 23125
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2248
timestamp 1626908933
transform 1 0 1200 0 1 23125
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1125
timestamp 1626908933
transform 1 0 1296 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3092
timestamp 1626908933
transform 1 0 1296 0 1 23643
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_672
timestamp 1626908933
transform 1 0 1440 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1394
timestamp 1626908933
transform 1 0 1440 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_568
timestamp 1626908933
transform 1 0 1056 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1166
timestamp 1626908933
transform 1 0 1056 0 -1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3138
timestamp 1626908933
transform 1 0 2448 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1171
timestamp 1626908933
transform 1 0 2448 0 1 23051
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1203
timestamp 1626908933
transform 1 0 2208 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_212
timestamp 1626908933
transform 1 0 2208 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1153
timestamp 1626908933
transform 1 0 2304 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_552
timestamp 1626908933
transform 1 0 2304 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_461
timestamp 1626908933
transform 1 0 2496 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_104
timestamp 1626908933
transform 1 0 2496 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3611
timestamp 1626908933
transform 1 0 2736 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1644
timestamp 1626908933
transform 1 0 2736 0 1 22977
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1154
timestamp 1626908933
transform 1 0 2592 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_553
timestamp 1626908933
transform 1 0 2592 0 -1 23976
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_942
timestamp 1626908933
transform 1 0 2900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_294
timestamp 1626908933
transform 1 0 2900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_942
timestamp 1626908933
transform 1 0 2900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_294
timestamp 1626908933
transform 1 0 2900 0 1 23310
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2257
timestamp 1626908933
transform 1 0 2928 0 1 23125
box -32 -32 32 32
use M1M2_PR  M1M2_PR_290
timestamp 1626908933
transform 1 0 2928 0 1 23125
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1915
timestamp 1626908933
transform 1 0 2784 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_924
timestamp 1626908933
transform 1 0 2784 0 -1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3660
timestamp 1626908933
transform 1 0 3024 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3128
timestamp 1626908933
transform 1 0 3120 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1725
timestamp 1626908933
transform 1 0 3024 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1193
timestamp 1626908933
transform 1 0 3120 0 1 23643
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_102
timestamp 1626908933
transform 1 0 2880 0 -1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_40
timestamp 1626908933
transform 1 0 2880 0 -1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_716
timestamp 1626908933
transform 1 0 3168 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_115
timestamp 1626908933
transform 1 0 3168 0 -1 23976
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1546
timestamp 1626908933
transform 1 0 3408 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3513
timestamp 1626908933
transform 1 0 3408 0 1 22977
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1636
timestamp 1626908933
transform 1 0 3408 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3571
timestamp 1626908933
transform 1 0 3408 0 1 22977
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_640
timestamp 1626908933
transform 1 0 3360 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1362
timestamp 1626908933
transform 1 0 3360 0 -1 23976
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1862
timestamp 1626908933
transform 1 0 3888 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3829
timestamp 1626908933
transform 1 0 3888 0 1 23199
box -32 -32 32 32
use L1M1_PR  L1M1_PR_310
timestamp 1626908933
transform 1 0 4368 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2245
timestamp 1626908933
transform 1 0 4368 0 1 22977
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1861
timestamp 1626908933
transform 1 0 3888 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3828
timestamp 1626908933
transform 1 0 3888 0 1 23643
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1836
timestamp 1626908933
transform 1 0 4272 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3771
timestamp 1626908933
transform 1 0 4272 0 1 23643
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_57
timestamp 1626908933
transform 1 0 4128 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_119
timestamp 1626908933
transform 1 0 4128 0 -1 23976
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2434
timestamp 1626908933
transform 1 0 4464 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_499
timestamp 1626908933
transform 1 0 4464 0 1 23421
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3837
timestamp 1626908933
transform 1 0 4560 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2255
timestamp 1626908933
transform 1 0 4464 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1870
timestamp 1626908933
transform 1 0 4560 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_288
timestamp 1626908933
transform 1 0 4464 0 1 22977
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1202
timestamp 1626908933
transform 1 0 4512 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_211
timestamp 1626908933
transform 1 0 4512 0 -1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3780
timestamp 1626908933
transform 1 0 4656 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3194
timestamp 1626908933
transform 1 0 4656 0 1 23199
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1845
timestamp 1626908933
transform 1 0 4656 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1259
timestamp 1626908933
transform 1 0 4656 0 1 23199
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2470
timestamp 1626908933
transform 1 0 4752 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_503
timestamp 1626908933
transform 1 0 4752 0 1 23421
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_270
timestamp 1626908933
transform 1 0 5300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_918
timestamp 1626908933
transform 1 0 5300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_270
timestamp 1626908933
transform 1 0 5300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_918
timestamp 1626908933
transform 1 0 5300 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_616
timestamp 1626908933
transform 1 0 4608 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1338
timestamp 1626908933
transform 1 0 4608 0 -1 23976
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3770
timestamp 1626908933
transform 1 0 5520 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1835
timestamp 1626908933
transform 1 0 5520 0 1 22977
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1100
timestamp 1626908933
transform 1 0 5376 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_502
timestamp 1626908933
transform 1 0 5376 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_210
timestamp 1626908933
transform 1 0 5760 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1201
timestamp 1626908933
transform 1 0 5760 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_518
timestamp 1626908933
transform 1 0 5808 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2485
timestamp 1626908933
transform 1 0 5808 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1855
timestamp 1626908933
transform 1 0 6096 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1856
timestamp 1626908933
transform 1 0 6000 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3822
timestamp 1626908933
transform 1 0 6096 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3823
timestamp 1626908933
transform 1 0 6000 0 1 23051
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_589
timestamp 1626908933
transform 1 0 5856 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1311
timestamp 1626908933
transform 1 0 5856 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_7
timestamp 1626908933
transform -1 0 7296 0 -1 23976
box -38 -49 710 715
use sky130_fd_sc_hs__a32oi_1  sky130_fd_sc_hs__a32oi_1_2
timestamp 1626908933
transform -1 0 7296 0 -1 23976
box -38 -49 710 715
use L1M1_PR  L1M1_PR_2366
timestamp 1626908933
transform 1 0 7152 0 1 23495
box -29 -23 29 23
use L1M1_PR  L1M1_PR_431
timestamp 1626908933
transform 1 0 7152 0 1 23495
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3164
timestamp 1626908933
transform 1 0 6960 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2401
timestamp 1626908933
transform 1 0 7152 0 1 23495
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1197
timestamp 1626908933
transform 1 0 6960 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_434
timestamp 1626908933
transform 1 0 7152 0 1 23495
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3766
timestamp 1626908933
transform 1 0 7344 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1831
timestamp 1626908933
transform 1 0 7344 0 1 23421
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_894
timestamp 1626908933
transform 1 0 7700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_246
timestamp 1626908933
transform 1 0 7700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_894
timestamp 1626908933
transform 1 0 7700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_246
timestamp 1626908933
transform 1 0 7700 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1200
timestamp 1626908933
transform 1 0 7584 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_209
timestamp 1626908933
transform 1 0 7584 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_460
timestamp 1626908933
transform 1 0 7488 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_103
timestamp 1626908933
transform 1 0 7488 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1155
timestamp 1626908933
transform 1 0 7296 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_554
timestamp 1626908933
transform 1 0 7296 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_553
timestamp 1626908933
transform 1 0 7680 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1275
timestamp 1626908933
transform 1 0 7680 0 -1 23976
box -38 -49 806 715
use L1M1_PR  L1M1_PR_513
timestamp 1626908933
transform 1 0 8400 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1249
timestamp 1626908933
transform 1 0 8688 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2448
timestamp 1626908933
transform 1 0 8400 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3184
timestamp 1626908933
transform 1 0 8688 0 1 23643
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_114
timestamp 1626908933
transform 1 0 8832 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_715
timestamp 1626908933
transform 1 0 8832 0 -1 23976
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1625
timestamp 1626908933
transform 1 0 9072 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3592
timestamp 1626908933
transform 1 0 9072 0 1 23051
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_534
timestamp 1626908933
transform 1 0 9024 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1256
timestamp 1626908933
transform 1 0 9024 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_53
timestamp 1626908933
transform -1 0 8832 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_115
timestamp 1626908933
transform -1 0 8832 0 -1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1091
timestamp 1626908933
transform 1 0 9840 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1095
timestamp 1626908933
transform 1 0 9264 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1186
timestamp 1626908933
transform 1 0 9456 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3058
timestamp 1626908933
transform 1 0 9840 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3062
timestamp 1626908933
transform 1 0 9264 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3153
timestamp 1626908933
transform 1 0 9456 0 1 23643
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1157
timestamp 1626908933
transform 1 0 9936 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3092
timestamp 1626908933
transform 1 0 9936 0 1 23421
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_34
timestamp 1626908933
transform -1 0 10368 0 -1 23976
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_73
timestamp 1626908933
transform -1 0 10368 0 -1 23976
box -38 -49 614 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_870
timestamp 1626908933
transform 1 0 10100 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_222
timestamp 1626908933
transform 1 0 10100 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_870
timestamp 1626908933
transform 1 0 10100 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_222
timestamp 1626908933
transform 1 0 10100 0 1 23310
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3096
timestamp 1626908933
transform 1 0 10128 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1161
timestamp 1626908933
transform 1 0 10128 0 1 23643
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2182
timestamp 1626908933
transform 1 0 10320 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_215
timestamp 1626908933
transform 1 0 10320 0 1 23643
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1199
timestamp 1626908933
transform 1 0 10368 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_208
timestamp 1626908933
transform 1 0 10368 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_509
timestamp 1626908933
transform 1 0 10464 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1231
timestamp 1626908933
transform 1 0 10464 0 -1 23976
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1006
timestamp 1626908933
transform 1 0 11088 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2973
timestamp 1626908933
transform 1 0 11088 0 1 23569
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1070
timestamp 1626908933
transform 1 0 11376 0 1 23569
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3005
timestamp 1626908933
transform 1 0 11376 0 1 23569
box -29 -23 29 23
use L1M1_PR  L1M1_PR_234
timestamp 1626908933
transform 1 0 11280 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2169
timestamp 1626908933
transform 1 0 11280 0 1 23643
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1009
timestamp 1626908933
transform 1 0 11664 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2976
timestamp 1626908933
transform 1 0 11664 0 1 23643
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1076
timestamp 1626908933
transform 1 0 11568 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3011
timestamp 1626908933
transform 1 0 11568 0 1 23643
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_65
timestamp 1626908933
transform -1 0 11808 0 -1 23976
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_26
timestamp 1626908933
transform -1 0 11808 0 -1 23976
box -38 -49 614 715
use L1M1_PR  L1M1_PR_3611
timestamp 1626908933
transform 1 0 11760 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1676
timestamp 1626908933
transform 1 0 11760 0 1 23421
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3553
timestamp 1626908933
transform 1 0 11856 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1586
timestamp 1626908933
transform 1 0 11856 0 1 23421
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1198
timestamp 1626908933
transform 1 0 12000 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_207
timestamp 1626908933
transform 1 0 12000 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_714
timestamp 1626908933
transform 1 0 11808 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_113
timestamp 1626908933
transform 1 0 11808 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_975
timestamp 1626908933
transform 1 0 12096 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_377
timestamp 1626908933
transform 1 0 12096 0 -1 23976
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_198
timestamp 1626908933
transform 1 0 12500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_846
timestamp 1626908933
transform 1 0 12500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_198
timestamp 1626908933
transform 1 0 12500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_846
timestamp 1626908933
transform 1 0 12500 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_102
timestamp 1626908933
transform 1 0 12480 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_459
timestamp 1626908933
transform 1 0 12480 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1614
timestamp 1626908933
transform 1 0 12720 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1615
timestamp 1626908933
transform 1 0 12720 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3581
timestamp 1626908933
transform 1 0 12720 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3582
timestamp 1626908933
transform 1 0 12720 0 1 23051
box -32 -32 32 32
use L1M1_PR  L1M1_PR_251
timestamp 1626908933
transform 1 0 13008 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2186
timestamp 1626908933
transform 1 0 13008 0 1 23421
box -29 -23 29 23
use M1M2_PR  M1M2_PR_229
timestamp 1626908933
transform 1 0 13296 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_230
timestamp 1626908933
transform 1 0 13296 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2196
timestamp 1626908933
transform 1 0 13296 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2197
timestamp 1626908933
transform 1 0 13296 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1721
timestamp 1626908933
transform 1 0 13488 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3688
timestamp 1626908933
transform 1 0 13488 0 1 23421
box -32 -32 32 32
use L1M1_PR  L1M1_PR_249
timestamp 1626908933
transform 1 0 13680 0 1 23199
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2184
timestamp 1626908933
transform 1 0 13680 0 1 23199
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_66
timestamp 1626908933
transform -1 0 15264 0 -1 23976
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_20
timestamp 1626908933
transform -1 0 15264 0 -1 23976
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1024
timestamp 1626908933
transform 1 0 13872 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2991
timestamp 1626908933
transform 1 0 13872 0 1 22977
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1092
timestamp 1626908933
transform 1 0 13872 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3027
timestamp 1626908933
transform 1 0 13872 0 1 22977
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1030
timestamp 1626908933
transform 1 0 14160 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2997
timestamp 1626908933
transform 1 0 14160 0 1 22977
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1098
timestamp 1626908933
transform 1 0 14064 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3033
timestamp 1626908933
transform 1 0 14064 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1668
timestamp 1626908933
transform 1 0 14256 0 1 23199
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3603
timestamp 1626908933
transform 1 0 14256 0 1 23199
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1608
timestamp 1626908933
transform 1 0 14640 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3575
timestamp 1626908933
transform 1 0 14640 0 1 23643
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1702
timestamp 1626908933
transform 1 0 14832 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3637
timestamp 1626908933
transform 1 0 14832 0 1 23643
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_174
timestamp 1626908933
transform 1 0 14900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_822
timestamp 1626908933
transform 1 0 14900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_174
timestamp 1626908933
transform 1 0 14900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_822
timestamp 1626908933
transform 1 0 14900 0 1 23310
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3546
timestamp 1626908933
transform 1 0 15216 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1579
timestamp 1626908933
transform 1 0 15216 0 1 23199
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3602
timestamp 1626908933
transform 1 0 15216 0 1 23569
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1667
timestamp 1626908933
transform 1 0 15216 0 1 23569
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3545
timestamp 1626908933
transform 1 0 15216 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1578
timestamp 1626908933
transform 1 0 15216 0 1 23569
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1197
timestamp 1626908933
transform 1 0 15456 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_206
timestamp 1626908933
transform 1 0 15456 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_713
timestamp 1626908933
transform 1 0 15264 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_112
timestamp 1626908933
transform 1 0 15264 0 -1 23976
box -38 -49 230 715
use M1M2_PR  M1M2_PR_240
timestamp 1626908933
transform 1 0 15504 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2207
timestamp 1626908933
transform 1 0 15504 0 1 23199
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2196
timestamp 1626908933
transform 1 0 15696 0 1 23199
box -29 -23 29 23
use L1M1_PR  L1M1_PR_261
timestamp 1626908933
transform 1 0 15696 0 1 23199
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3012
timestamp 1626908933
transform 1 0 15696 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1045
timestamp 1626908933
transform 1 0 15696 0 1 23643
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1196
timestamp 1626908933
transform 1 0 16320 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_205
timestamp 1626908933
transform 1 0 16320 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1126
timestamp 1626908933
transform 1 0 15552 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_404
timestamp 1626908933
transform 1 0 15552 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1156
timestamp 1626908933
transform 1 0 16416 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_555
timestamp 1626908933
transform 1 0 16416 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_204
timestamp 1626908933
transform 1 0 16992 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1195
timestamp 1626908933
transform 1 0 16992 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1708
timestamp 1626908933
transform 1 0 16656 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3675
timestamp 1626908933
transform 1 0 16656 0 1 23051
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1111
timestamp 1626908933
transform 1 0 16752 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1662
timestamp 1626908933
transform 1 0 16944 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3046
timestamp 1626908933
transform 1 0 16752 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3597
timestamp 1626908933
transform 1 0 16944 0 1 23421
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_150
timestamp 1626908933
transform 1 0 17300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_798
timestamp 1626908933
transform 1 0 17300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_150
timestamp 1626908933
transform 1 0 17300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_798
timestamp 1626908933
transform 1 0 17300 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_279
timestamp 1626908933
transform 1 0 17088 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_877
timestamp 1626908933
transform 1 0 17088 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_43
timestamp 1626908933
transform 1 0 16608 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_105
timestamp 1626908933
transform 1 0 16608 0 -1 23976
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3632
timestamp 1626908933
transform 1 0 17520 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1697
timestamp 1626908933
transform 1 0 17520 0 1 22977
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3570
timestamp 1626908933
transform 1 0 17520 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1603
timestamp 1626908933
transform 1 0 17520 0 1 22977
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1194
timestamp 1626908933
transform 1 0 17568 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_203
timestamp 1626908933
transform 1 0 17568 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_458
timestamp 1626908933
transform 1 0 17472 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_101
timestamp 1626908933
transform 1 0 17472 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3540
timestamp 1626908933
transform 1 0 17808 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3539
timestamp 1626908933
transform 1 0 17808 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1573
timestamp 1626908933
transform 1 0 17808 0 1 23051
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1572
timestamp 1626908933
transform 1 0 17808 0 1 23421
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_202
timestamp 1626908933
transform 1 0 18048 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1193
timestamp 1626908933
transform 1 0 18048 0 -1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1661
timestamp 1626908933
transform 1 0 17904 0 1 23051
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3596
timestamp 1626908933
transform 1 0 17904 0 1 23051
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_351
timestamp 1626908933
transform 1 0 18144 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1073
timestamp 1626908933
transform 1 0 18144 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_264
timestamp 1626908933
transform 1 0 17664 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_862
timestamp 1626908933
transform 1 0 17664 0 -1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3275
timestamp 1626908933
transform 1 0 18960 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1308
timestamp 1626908933
transform 1 0 18960 0 1 22977
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1192
timestamp 1626908933
transform 1 0 18912 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_201
timestamp 1626908933
transform 1 0 18912 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_835
timestamp 1626908933
transform 1 0 19008 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_237
timestamp 1626908933
transform 1 0 19008 0 -1 23976
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3323
timestamp 1626908933
transform 1 0 19152 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1388
timestamp 1626908933
transform 1 0 19152 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1380
timestamp 1626908933
transform 1 0 19536 0 1 23125
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3315
timestamp 1626908933
transform 1 0 19536 0 1 23125
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_126
timestamp 1626908933
transform 1 0 19700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_774
timestamp 1626908933
transform 1 0 19700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_126
timestamp 1626908933
transform 1 0 19700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_774
timestamp 1626908933
transform 1 0 19700 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_200
timestamp 1626908933
transform 1 0 20160 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1191
timestamp 1626908933
transform 1 0 20160 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_324
timestamp 1626908933
transform 1 0 19392 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1046
timestamp 1626908933
transform 1 0 19392 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_813
timestamp 1626908933
transform 1 0 20256 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_215
timestamp 1626908933
transform 1 0 20256 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1018
timestamp 1626908933
transform 1 0 20640 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_296
timestamp 1626908933
transform 1 0 20640 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1190
timestamp 1626908933
transform 1 0 21600 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_199
timestamp 1626908933
transform 1 0 21600 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_712
timestamp 1626908933
transform 1 0 21408 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_111
timestamp 1626908933
transform 1 0 21408 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_990
timestamp 1626908933
transform 1 0 21696 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_268
timestamp 1626908933
transform 1 0 21696 0 -1 23976
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_750
timestamp 1626908933
transform 1 0 22100 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_102
timestamp 1626908933
transform 1 0 22100 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_750
timestamp 1626908933
transform 1 0 22100 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_102
timestamp 1626908933
transform 1 0 22100 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_100
timestamp 1626908933
transform 1 0 22464 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_457
timestamp 1626908933
transform 1 0 22464 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_421
timestamp 1626908933
transform 1 0 22608 0 1 23199
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2388
timestamp 1626908933
transform 1 0 22608 0 1 23199
box -32 -32 32 32
use L1M1_PR  L1M1_PR_417
timestamp 1626908933
transform 1 0 22608 0 1 23199
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1513
timestamp 1626908933
transform 1 0 22800 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2352
timestamp 1626908933
transform 1 0 22608 0 1 23199
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3448
timestamp 1626908933
transform 1 0 22800 0 1 22977
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_245
timestamp 1626908933
transform 1 0 22560 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_967
timestamp 1626908933
transform 1 0 22560 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_711
timestamp 1626908933
transform 1 0 23328 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_110
timestamp 1626908933
transform 1 0 23328 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_754
timestamp 1626908933
transform 1 0 23520 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_156
timestamp 1626908933
transform 1 0 23520 0 -1 23976
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3756
timestamp 1626908933
transform 1 0 24144 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1821
timestamp 1626908933
transform 1 0 24144 0 1 22977
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3807
timestamp 1626908933
transform 1 0 24144 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1840
timestamp 1626908933
transform 1 0 24144 0 1 22977
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2348
timestamp 1626908933
transform 1 0 24336 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_413
timestamp 1626908933
transform 1 0 24336 0 1 22977
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2385
timestamp 1626908933
transform 1 0 24240 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_418
timestamp 1626908933
transform 1 0 24240 0 1 22977
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3801
timestamp 1626908933
transform 1 0 24432 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1866
timestamp 1626908933
transform 1 0 24432 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3737
timestamp 1626908933
transform 1 0 24624 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1802
timestamp 1626908933
transform 1 0 24624 0 1 22977
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_726
timestamp 1626908933
transform 1 0 24500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_78
timestamp 1626908933
transform 1 0 24500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_726
timestamp 1626908933
transform 1 0 24500 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_78
timestamp 1626908933
transform 1 0 24500 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_215
timestamp 1626908933
transform 1 0 23904 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_937
timestamp 1626908933
transform 1 0 23904 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1189
timestamp 1626908933
transform 1 0 24672 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_198
timestamp 1626908933
transform 1 0 24672 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_729
timestamp 1626908933
transform 1 0 24768 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_131
timestamp 1626908933
transform 1 0 24768 0 -1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3375
timestamp 1626908933
transform 1 0 25392 0 1 23125
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3255
timestamp 1626908933
transform 1 0 25200 0 1 23125
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1408
timestamp 1626908933
transform 1 0 25392 0 1 23125
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1288
timestamp 1626908933
transform 1 0 25200 0 1 23125
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_902
timestamp 1626908933
transform 1 0 25152 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_180
timestamp 1626908933
transform 1 0 25152 0 -1 23976
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3426
timestamp 1626908933
transform 1 0 26352 0 1 23125
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1491
timestamp 1626908933
transform 1 0 26352 0 1 23125
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_710
timestamp 1626908933
transform 1 0 25920 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_109
timestamp 1626908933
transform 1 0 25920 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_701
timestamp 1626908933
transform 1 0 26112 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_103
timestamp 1626908933
transform 1 0 26112 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_873
timestamp 1626908933
transform 1 0 26496 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_151
timestamp 1626908933
transform 1 0 26496 0 -1 23976
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_54
timestamp 1626908933
transform 1 0 26900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_702
timestamp 1626908933
transform 1 0 26900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_54
timestamp 1626908933
transform 1 0 26900 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_702
timestamp 1626908933
transform 1 0 26900 0 1 23310
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1775
timestamp 1626908933
transform 1 0 27120 0 1 23125
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3742
timestamp 1626908933
transform 1 0 27120 0 1 23125
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_197
timestamp 1626908933
transform 1 0 27264 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_925
timestamp 1626908933
transform 1 0 27360 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1188
timestamp 1626908933
transform 1 0 27264 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1916
timestamp 1626908933
transform 1 0 27360 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3774
timestamp 1626908933
transform 1 0 27504 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1807
timestamp 1626908933
transform 1 0 27504 0 1 22977
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_709
timestamp 1626908933
transform 1 0 27552 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_108
timestamp 1626908933
transform 1 0 27552 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_456
timestamp 1626908933
transform 1 0 27456 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_99
timestamp 1626908933
transform 1 0 27456 0 -1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_415
timestamp 1626908933
transform 1 0 27888 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1892
timestamp 1626908933
transform 1 0 28368 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2382
timestamp 1626908933
transform 1 0 27888 0 1 22977
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3859
timestamp 1626908933
transform 1 0 28368 0 1 22977
box -32 -32 32 32
use L1M1_PR  L1M1_PR_411
timestamp 1626908933
transform 1 0 28272 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1864
timestamp 1626908933
transform 1 0 28368 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2346
timestamp 1626908933
transform 1 0 28272 0 1 22977
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3799
timestamp 1626908933
transform 1 0 28368 0 1 22977
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_120
timestamp 1626908933
transform 1 0 27744 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_842
timestamp 1626908933
transform 1 0 27744 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_196
timestamp 1626908933
transform 1 0 28896 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1187
timestamp 1626908933
transform 1 0 28896 0 -1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1791
timestamp 1626908933
transform 1 0 28560 0 1 23125
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3726
timestamp 1626908933
transform 1 0 28560 0 1 23125
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1888
timestamp 1626908933
transform 1 0 29040 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3855
timestamp 1626908933
transform 1 0 29040 0 1 23569
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_30
timestamp 1626908933
transform 1 0 29300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_678
timestamp 1626908933
transform 1 0 29300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_30
timestamp 1626908933
transform 1 0 29300 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_678
timestamp 1626908933
transform 1 0 29300 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_86
timestamp 1626908933
transform 1 0 28992 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_808
timestamp 1626908933
transform 1 0 28992 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_59
timestamp 1626908933
transform 1 0 28512 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_657
timestamp 1626908933
transform 1 0 28512 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_25
timestamp 1626908933
transform 1 0 30144 0 -1 23976
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_10
timestamp 1626908933
transform 1 0 30144 0 -1 23976
box -38 -49 710 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_626
timestamp 1626908933
transform 1 0 29760 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_28
timestamp 1626908933
transform 1 0 29760 0 -1 23976
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3746
timestamp 1626908933
transform 1 0 30192 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1811
timestamp 1626908933
transform 1 0 30192 0 1 23643
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3854
timestamp 1626908933
transform 1 0 30288 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3745
timestamp 1626908933
transform 1 0 30288 0 1 23421
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1887
timestamp 1626908933
transform 1 0 30288 0 1 23569
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1778
timestamp 1626908933
transform 1 0 30288 0 1 23421
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3794
timestamp 1626908933
transform 1 0 30576 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2341
timestamp 1626908933
transform 1 0 30480 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1859
timestamp 1626908933
transform 1 0 30576 0 1 23643
box -29 -23 29 23
use L1M1_PR  L1M1_PR_406
timestamp 1626908933
transform 1 0 30480 0 1 23643
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2379
timestamp 1626908933
transform 1 0 30480 0 1 23643
box -32 -32 32 32
use M1M2_PR  M1M2_PR_412
timestamp 1626908933
transform 1 0 30480 0 1 23643
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3727
timestamp 1626908933
transform 1 0 30768 0 1 23421
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1792
timestamp 1626908933
transform 1 0 30768 0 1 23421
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1186
timestamp 1626908933
transform 1 0 30816 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_195
timestamp 1626908933
transform 1 0 30816 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_25
timestamp 1626908933
transform 1 0 30912 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_747
timestamp 1626908933
transform 1 0 30912 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_98
timestamp 1626908933
transform 1 0 31680 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_455
timestamp 1626908933
transform 1 0 31680 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_556
timestamp 1626908933
transform 1 0 31776 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1157
timestamp 1626908933
transform 1 0 31776 0 -1 23976
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_6
timestamp 1626908933
transform 1 0 31700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_654
timestamp 1626908933
transform 1 0 31700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_6
timestamp 1626908933
transform 1 0 31700 0 1 23310
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_654
timestamp 1626908933
transform 1 0 31700 0 1 23310
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_926
timestamp 1626908933
transform 1 0 31968 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1917
timestamp 1626908933
transform 1 0 31968 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_97
timestamp 1626908933
transform 1 0 288 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_454
timestamp 1626908933
transform 1 0 288 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_557
timestamp 1626908933
transform 1 0 0 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1158
timestamp 1626908933
transform 1 0 0 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_194
timestamp 1626908933
transform 1 0 384 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_927
timestamp 1626908933
transform 1 0 192 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1185
timestamp 1626908933
transform 1 0 384 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1918
timestamp 1626908933
transform 1 0 192 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_693
timestamp 1626908933
transform 1 0 480 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1415
timestamp 1626908933
transform 1 0 480 0 1 23976
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1128
timestamp 1626908933
transform 1 0 1488 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3095
timestamp 1626908933
transform 1 0 1488 0 1 23865
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_630
timestamp 1626908933
transform 1 0 1700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1278
timestamp 1626908933
transform 1 0 1700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_630
timestamp 1626908933
transform 1 0 1700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1278
timestamp 1626908933
transform 1 0 1700 0 1 23976
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3131
timestamp 1626908933
transform 1 0 1296 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1196
timestamp 1626908933
transform 1 0 1296 0 1 24235
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3091
timestamp 1626908933
transform 1 0 1296 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1124
timestamp 1626908933
transform 1 0 1296 0 1 24235
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3137
timestamp 1626908933
transform 1 0 1680 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1202
timestamp 1626908933
transform 1 0 1680 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3134
timestamp 1626908933
transform 1 0 1392 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1199
timestamp 1626908933
transform 1 0 1392 0 1 24309
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3094
timestamp 1626908933
transform 1 0 1680 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1127
timestamp 1626908933
transform 1 0 1680 0 1 24309
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_4
timestamp 1626908933
transform 1 0 1632 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_56
timestamp 1626908933
transform 1 0 1632 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_51
timestamp 1626908933
transform 1 0 1248 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_113
timestamp 1626908933
transform 1 0 1248 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1184
timestamp 1626908933
transform 1 0 2016 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_193
timestamp 1626908933
transform 1 0 2016 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1382
timestamp 1626908933
transform 1 0 2112 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_660
timestamp 1626908933
transform 1 0 2112 0 1 23976
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3133
timestamp 1626908933
transform 1 0 2832 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1198
timestamp 1626908933
transform 1 0 2832 0 1 23865
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3098
timestamp 1626908933
transform 1 0 2928 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3097
timestamp 1626908933
transform 1 0 2928 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1131
timestamp 1626908933
transform 1 0 2928 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1130
timestamp 1626908933
transform 1 0 2928 0 1 24087
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1183
timestamp 1626908933
transform 1 0 2880 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_192
timestamp 1626908933
transform 1 0 2880 0 1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3135
timestamp 1626908933
transform 1 0 3024 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1200
timestamp 1626908933
transform 1 0 3024 0 1 23865
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_639
timestamp 1626908933
transform 1 0 3360 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1361
timestamp 1626908933
transform 1 0 3360 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_542
timestamp 1626908933
transform 1 0 2976 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1140
timestamp 1626908933
transform 1 0 2976 0 1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1205
timestamp 1626908933
transform 1 0 4368 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3172
timestamp 1626908933
transform 1 0 4368 0 1 23717
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1273
timestamp 1626908933
transform 1 0 4176 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3208
timestamp 1626908933
transform 1 0 4176 0 1 23717
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_606
timestamp 1626908933
transform 1 0 4100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1254
timestamp 1626908933
transform 1 0 4100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_606
timestamp 1626908933
transform 1 0 4100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1254
timestamp 1626908933
transform 1 0 4100 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1204
timestamp 1626908933
transform 1 0 4368 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3171
timestamp 1626908933
transform 1 0 4368 0 1 24087
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1272
timestamp 1626908933
transform 1 0 4272 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1283
timestamp 1626908933
transform 1 0 4368 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1846
timestamp 1626908933
transform 1 0 4176 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3207
timestamp 1626908933
transform 1 0 4272 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3218
timestamp 1626908933
transform 1 0 4368 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3781
timestamp 1626908933
transform 1 0 4176 0 1 24235
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_59
timestamp 1626908933
transform -1 0 4512 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_121
timestamp 1626908933
transform -1 0 4512 0 1 23976
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1275
timestamp 1626908933
transform 1 0 4464 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3210
timestamp 1626908933
transform 1 0 4464 0 1 23717
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1213
timestamp 1626908933
transform 1 0 4464 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1869
timestamp 1626908933
transform 1 0 4560 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3180
timestamp 1626908933
transform 1 0 4464 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3836
timestamp 1626908933
transform 1 0 4560 0 1 24161
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1285
timestamp 1626908933
transform 1 0 4464 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3220
timestamp 1626908933
transform 1 0 4464 0 1 24235
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_191
timestamp 1626908933
transform 1 0 4512 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1182
timestamp 1626908933
transform 1 0 4512 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_96
timestamp 1626908933
transform 1 0 4992 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_453
timestamp 1626908933
transform 1 0 4992 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_107
timestamp 1626908933
transform 1 0 5088 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_708
timestamp 1626908933
transform 1 0 5088 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_501
timestamp 1626908933
transform 1 0 5280 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_515
timestamp 1626908933
transform 1 0 4608 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1099
timestamp 1626908933
transform 1 0 5280 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1113
timestamp 1626908933
transform 1 0 4608 0 1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3174
timestamp 1626908933
transform 1 0 5808 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2478
timestamp 1626908933
transform 1 0 5712 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1207
timestamp 1626908933
transform 1 0 5808 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_511
timestamp 1626908933
transform 1 0 5712 0 1 23865
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3775
timestamp 1626908933
transform 1 0 5904 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2442
timestamp 1626908933
transform 1 0 5712 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1840
timestamp 1626908933
transform 1 0 5904 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_507
timestamp 1626908933
transform 1 0 5712 0 1 24235
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2479
timestamp 1626908933
transform 1 0 5616 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_512
timestamp 1626908933
transform 1 0 5616 0 1 24235
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_114
timestamp 1626908933
transform 1 0 5664 0 1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_53
timestamp 1626908933
transform 1 0 5664 0 1 23976
box -38 -49 326 715
use M1M2_PR  M1M2_PR_516
timestamp 1626908933
transform 1 0 6288 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2483
timestamp 1626908933
transform 1 0 6288 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1864
timestamp 1626908933
transform 1 0 6768 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3831
timestamp 1626908933
transform 1 0 6768 0 1 23717
box -32 -32 32 32
use L1M1_PR  L1M1_PR_511
timestamp 1626908933
transform 1 0 6672 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2446
timestamp 1626908933
transform 1 0 6672 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_506
timestamp 1626908933
transform 1 0 6864 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2441
timestamp 1626908933
transform 1 0 6864 0 1 23865
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_582
timestamp 1626908933
transform 1 0 6500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1230
timestamp 1626908933
transform 1 0 6500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_582
timestamp 1626908933
transform 1 0 6500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1230
timestamp 1626908933
transform 1 0 6500 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3833
timestamp 1626908933
transform 1 0 6672 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3178
timestamp 1626908933
transform 1 0 6672 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1866
timestamp 1626908933
transform 1 0 6672 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1211
timestamp 1626908933
transform 1 0 6672 0 1 24309
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_0
timestamp 1626908933
transform 1 0 6720 0 1 23976
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_8
timestamp 1626908933
transform 1 0 6720 0 1 23976
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_588
timestamp 1626908933
transform 1 0 5952 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1310
timestamp 1626908933
transform 1 0 5952 0 1 23976
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3773
timestamp 1626908933
transform 1 0 6960 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2449
timestamp 1626908933
transform 1 0 7056 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1838
timestamp 1626908933
transform 1 0 6960 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_514
timestamp 1626908933
transform 1 0 7056 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3193
timestamp 1626908933
transform 1 0 6960 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3192
timestamp 1626908933
transform 1 0 7056 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1258
timestamp 1626908933
transform 1 0 6960 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1257
timestamp 1626908933
transform 1 0 7056 0 1 24309
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3163
timestamp 1626908933
transform 1 0 6960 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1196
timestamp 1626908933
transform 1 0 6960 0 1 24309
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_928
timestamp 1626908933
transform 1 0 7200 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1919
timestamp 1626908933
transform 1 0 7200 0 1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_296
timestamp 1626908933
transform 1 0 7632 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2231
timestamp 1626908933
transform 1 0 7632 0 1 24087
box -29 -23 29 23
use M1M2_PR  M1M2_PR_272
timestamp 1626908933
transform 1 0 7920 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_273
timestamp 1626908933
transform 1 0 7920 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1741
timestamp 1626908933
transform 1 0 7920 0 1 24457
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2239
timestamp 1626908933
transform 1 0 7920 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2240
timestamp 1626908933
transform 1 0 7920 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3708
timestamp 1626908933
transform 1 0 7920 0 1 24457
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_69
timestamp 1626908933
transform -1 0 9984 0 1 23976
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_23
timestamp 1626908933
transform -1 0 9984 0 1 23976
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1191
timestamp 1626908933
transform 1 0 8304 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3158
timestamp 1626908933
transform 1 0 8304 0 1 23717
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1252
timestamp 1626908933
transform 1 0 8496 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3187
timestamp 1626908933
transform 1 0 8496 0 1 23717
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1188
timestamp 1626908933
transform 1 0 8784 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3155
timestamp 1626908933
transform 1 0 8784 0 1 23717
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1250
timestamp 1626908933
transform 1 0 8784 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3185
timestamp 1626908933
transform 1 0 8784 0 1 23717
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_558
timestamp 1626908933
transform 1 0 8900 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1206
timestamp 1626908933
transform 1 0 8900 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_558
timestamp 1626908933
transform 1 0 8900 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1206
timestamp 1626908933
transform 1 0 8900 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1628
timestamp 1626908933
transform 1 0 8688 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3595
timestamp 1626908933
transform 1 0 8688 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1624
timestamp 1626908933
transform 1 0 9072 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3591
timestamp 1626908933
transform 1 0 9072 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1195
timestamp 1626908933
transform 1 0 9456 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3162
timestamp 1626908933
transform 1 0 9456 0 1 24309
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1712
timestamp 1626908933
transform 1 0 9552 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3647
timestamp 1626908933
transform 1 0 9552 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_293
timestamp 1626908933
transform 1 0 9744 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2228
timestamp 1626908933
transform 1 0 9744 0 1 23865
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_95
timestamp 1626908933
transform 1 0 9984 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_452
timestamp 1626908933
transform 1 0 9984 0 1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1644
timestamp 1626908933
transform 1 0 9936 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3579
timestamp 1626908933
transform 1 0 9936 0 1 24235
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1555
timestamp 1626908933
transform 1 0 10128 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3522
timestamp 1626908933
transform 1 0 10128 0 1 23865
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1643
timestamp 1626908933
transform 1 0 10320 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3578
timestamp 1626908933
transform 1 0 10320 0 1 23865
box -29 -23 29 23
use M1M2_PR  M1M2_PR_214
timestamp 1626908933
transform 1 0 10320 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_242
timestamp 1626908933
transform 1 0 10608 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1554
timestamp 1626908933
transform 1 0 10128 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2181
timestamp 1626908933
transform 1 0 10320 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2209
timestamp 1626908933
transform 1 0 10608 0 1 24235
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3521
timestamp 1626908933
transform 1 0 10128 0 1 24235
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_508
timestamp 1626908933
transform 1 0 10464 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1230
timestamp 1626908933
transform 1 0 10464 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_418
timestamp 1626908933
transform 1 0 10080 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1016
timestamp 1626908933
transform 1 0 10080 0 1 23976
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_534
timestamp 1626908933
transform 1 0 11300 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1182
timestamp 1626908933
transform 1 0 11300 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_534
timestamp 1626908933
transform 1 0 11300 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1182
timestamp 1626908933
transform 1 0 11300 0 1 23976
box -100 -49 100 49
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_48
timestamp 1626908933
transform 1 0 11616 0 1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_109
timestamp 1626908933
transform 1 0 11616 0 1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_106
timestamp 1626908933
transform 1 0 11904 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_707
timestamp 1626908933
transform 1 0 11904 0 1 23976
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1008
timestamp 1626908933
transform 1 0 11664 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2975
timestamp 1626908933
transform 1 0 11664 0 1 24161
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1074
timestamp 1626908933
transform 1 0 11760 0 1 24161
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3009
timestamp 1626908933
transform 1 0 11760 0 1 24161
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_3
timestamp 1626908933
transform 1 0 11232 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_55
timestamp 1626908933
transform 1 0 11232 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_190
timestamp 1626908933
transform 1 0 12096 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1181
timestamp 1626908933
transform 1 0 12096 0 1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_232
timestamp 1626908933
transform 1 0 12048 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2199
timestamp 1626908933
transform 1 0 12048 0 1 23865
box -32 -32 32 32
use L1M1_PR  L1M1_PR_233
timestamp 1626908933
transform 1 0 11952 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2168
timestamp 1626908933
transform 1 0 11952 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_252
timestamp 1626908933
transform 1 0 12720 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2187
timestamp 1626908933
transform 1 0 12720 0 1 23865
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_469
timestamp 1626908933
transform 1 0 12192 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1191
timestamp 1626908933
transform 1 0 12192 0 1 23976
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2189
timestamp 1626908933
transform 1 0 13008 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_254
timestamp 1626908933
transform 1 0 13008 0 1 24309
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2201
timestamp 1626908933
transform 1 0 13008 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_234
timestamp 1626908933
transform 1 0 13008 0 1 24309
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1160
timestamp 1626908933
transform 1 0 13440 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_438
timestamp 1626908933
transform 1 0 13440 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_45
timestamp 1626908933
transform 1 0 12960 0 1 23976
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_114
timestamp 1626908933
transform 1 0 12960 0 1 23976
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1158
timestamp 1626908933
transform 1 0 13700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_510
timestamp 1626908933
transform 1 0 13700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1158
timestamp 1626908933
transform 1 0 13700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_510
timestamp 1626908933
transform 1 0 13700 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1029
timestamp 1626908933
transform 1 0 14160 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2996
timestamp 1626908933
transform 1 0 14160 0 1 24309
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_49
timestamp 1626908933
transform -1 0 14496 0 1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_111
timestamp 1626908933
transform -1 0 14496 0 1 23976
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_189
timestamp 1626908933
transform 1 0 14496 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1180
timestamp 1626908933
transform 1 0 14496 0 1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1033
timestamp 1626908933
transform 1 0 14352 0 1 24457
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3000
timestamp 1626908933
transform 1 0 14352 0 1 24457
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1095
timestamp 1626908933
transform 1 0 14256 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3030
timestamp 1626908933
transform 1 0 14256 0 1 24309
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_331
timestamp 1626908933
transform 1 0 14592 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_929
timestamp 1626908933
transform 1 0 14592 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_94
timestamp 1626908933
transform 1 0 14976 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_451
timestamp 1626908933
transform 1 0 14976 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_558
timestamp 1626908933
transform 1 0 15072 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1159
timestamp 1626908933
transform 1 0 15072 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_929
timestamp 1626908933
transform 1 0 15264 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1920
timestamp 1626908933
transform 1 0 15264 0 1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_239
timestamp 1626908933
transform 1 0 15504 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2206
timestamp 1626908933
transform 1 0 15504 0 1 24309
box -32 -32 32 32
use L1M1_PR  L1M1_PR_262
timestamp 1626908933
transform 1 0 15504 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2197
timestamp 1626908933
transform 1 0 15504 0 1 24309
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_115
timestamp 1626908933
transform -1 0 15840 0 1 23976
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_46
timestamp 1626908933
transform -1 0 15840 0 1 23976
box -38 -49 518 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_486
timestamp 1626908933
transform 1 0 16100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1134
timestamp 1626908933
transform 1 0 16100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_486
timestamp 1626908933
transform 1 0 16100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1134
timestamp 1626908933
transform 1 0 16100 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1044
timestamp 1626908933
transform 1 0 15696 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3011
timestamp 1626908933
transform 1 0 15696 0 1 24087
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1112
timestamp 1626908933
transform 1 0 15696 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3047
timestamp 1626908933
transform 1 0 15696 0 1 24087
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_390
timestamp 1626908933
transform 1 0 16224 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1112
timestamp 1626908933
transform 1 0 16224 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_301
timestamp 1626908933
transform 1 0 15840 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_899
timestamp 1626908933
transform 1 0 15840 0 1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3009
timestamp 1626908933
transform 1 0 16464 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1042
timestamp 1626908933
transform 1 0 16464 0 1 23717
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_188
timestamp 1626908933
transform 1 0 16992 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1179
timestamp 1626908933
transform 1 0 16992 0 1 23976
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1047
timestamp 1626908933
transform 1 0 16848 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3014
timestamp 1626908933
transform 1 0 16848 0 1 23717
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1106
timestamp 1626908933
transform 1 0 16656 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1113
timestamp 1626908933
transform 1 0 16944 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3041
timestamp 1626908933
transform 1 0 16656 0 1 23717
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3048
timestamp 1626908933
transform 1 0 16944 0 1 23717
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_278
timestamp 1626908933
transform 1 0 17088 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_876
timestamp 1626908933
transform 1 0 17088 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1178
timestamp 1626908933
transform 1 0 18240 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_187
timestamp 1626908933
transform 1 0 18240 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1088
timestamp 1626908933
transform 1 0 17472 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_366
timestamp 1626908933
transform 1 0 17472 0 1 23976
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_462
timestamp 1626908933
transform 1 0 18500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1110
timestamp 1626908933
transform 1 0 18500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_462
timestamp 1626908933
transform 1 0 18500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1110
timestamp 1626908933
transform 1 0 18500 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1307
timestamp 1626908933
transform 1 0 18960 0 1 24457
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3274
timestamp 1626908933
transform 1 0 18960 0 1 24457
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_336
timestamp 1626908933
transform 1 0 18720 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1058
timestamp 1626908933
transform 1 0 18720 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_248
timestamp 1626908933
transform 1 0 18336 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_846
timestamp 1626908933
transform 1 0 18336 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_228
timestamp 1626908933
transform 1 0 19488 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_826
timestamp 1626908933
transform 1 0 19488 0 1 23976
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2302
timestamp 1626908933
transform 1 0 19920 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_335
timestamp 1626908933
transform 1 0 19920 0 1 24309
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1921
timestamp 1626908933
transform 1 0 19872 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_930
timestamp 1626908933
transform 1 0 19872 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_450
timestamp 1626908933
transform 1 0 19968 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_93
timestamp 1626908933
transform 1 0 19968 0 1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3379
timestamp 1626908933
transform 1 0 20208 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1444
timestamp 1626908933
transform 1 0 20208 0 1 24087
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3327
timestamp 1626908933
transform 1 0 20208 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1360
timestamp 1626908933
transform 1 0 20208 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1286
timestamp 1626908933
transform 1 0 20400 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3253
timestamp 1626908933
transform 1 0 20400 0 1 24383
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1379
timestamp 1626908933
transform 1 0 20400 0 1 24383
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3314
timestamp 1626908933
transform 1 0 20400 0 1 24383
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1294
timestamp 1626908933
transform 1 0 21168 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3261
timestamp 1626908933
transform 1 0 21168 0 1 24383
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1383
timestamp 1626908933
transform 1 0 21168 0 1 24383
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3318
timestamp 1626908933
transform 1 0 21168 0 1 24383
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_438
timestamp 1626908933
transform 1 0 20900 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1086
timestamp 1626908933
transform 1 0 20900 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_438
timestamp 1626908933
transform 1 0 20900 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1086
timestamp 1626908933
transform 1 0 20900 0 1 23976
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1383
timestamp 1626908933
transform 1 0 21648 0 1 24161
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3350
timestamp 1626908933
transform 1 0 21648 0 1 24161
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_183
timestamp 1626908933
transform 1 0 22080 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_781
timestamp 1626908933
transform 1 0 22080 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_105
timestamp 1626908933
transform 1 0 21888 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_706
timestamp 1626908933
transform 1 0 21888 0 1 23976
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1386
timestamp 1626908933
transform 1 0 21744 0 1 24383
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3321
timestamp 1626908933
transform 1 0 21744 0 1 24383
box -29 -23 29 23
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_23
timestamp 1626908933
transform -1 0 21888 0 1 23976
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_11
timestamp 1626908933
transform -1 0 21888 0 1 23976
box -38 -49 1862 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_414
timestamp 1626908933
transform 1 0 23300 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1062
timestamp 1626908933
transform 1 0 23300 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_414
timestamp 1626908933
transform 1 0 23300 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1062
timestamp 1626908933
transform 1 0 23300 0 1 23976
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1463
timestamp 1626908933
transform 1 0 22800 0 1 24235
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3398
timestamp 1626908933
transform 1 0 22800 0 1 24235
box -29 -23 29 23
use M1M2_PR  M1M2_PR_420
timestamp 1626908933
transform 1 0 22608 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2387
timestamp 1626908933
transform 1 0 22608 0 1 24309
box -32 -32 32 32
use L1M1_PR  L1M1_PR_416
timestamp 1626908933
transform 1 0 22608 0 1 24309
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2351
timestamp 1626908933
transform 1 0 22608 0 1 24309
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1301
timestamp 1626908933
transform 1 0 23472 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3268
timestamp 1626908933
transform 1 0 23472 0 1 24383
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2329
timestamp 1626908933
transform 1 0 24720 0 1 24087
box -29 -23 29 23
use L1M1_PR  L1M1_PR_394
timestamp 1626908933
transform 1 0 24720 0 1 24087
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2355
timestamp 1626908933
transform 1 0 23664 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2338
timestamp 1626908933
transform 1 0 24336 0 1 24087
box -32 -32 32 32
use M1M2_PR  M1M2_PR_388
timestamp 1626908933
transform 1 0 23664 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_371
timestamp 1626908933
transform 1 0 24336 0 1 24087
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1922
timestamp 1626908933
transform 1 0 24864 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_931
timestamp 1626908933
transform 1 0 24864 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_5
timestamp 1626908933
transform 1 0 22464 0 1 23976
box -38 -49 2438 715
use sky130_fd_sc_hs__dfstp_2  sky130_fd_sc_hs__dfstp_2_1
timestamp 1626908933
transform 1 0 22464 0 1 23976
box -38 -49 2438 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_92
timestamp 1626908933
transform 1 0 24960 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_449
timestamp 1626908933
transform 1 0 24960 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_122
timestamp 1626908933
transform 1 0 25152 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_720
timestamp 1626908933
transform 1 0 25152 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_186
timestamp 1626908933
transform 1 0 25056 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1177
timestamp 1626908933
transform 1 0 25056 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_185
timestamp 1626908933
transform 1 0 25536 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1176
timestamp 1626908933
transform 1 0 25536 0 1 23976
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_390
timestamp 1626908933
transform 1 0 25700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1038
timestamp 1626908933
transform 1 0 25700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_390
timestamp 1626908933
transform 1 0 25700 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1038
timestamp 1626908933
transform 1 0 25700 0 1 23976
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1371
timestamp 1626908933
transform 1 0 25968 0 1 24383
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3306
timestamp 1626908933
transform 1 0 25968 0 1 24383
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1279
timestamp 1626908933
transform 1 0 26352 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3246
timestamp 1626908933
transform 1 0 26352 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1298
timestamp 1626908933
transform 1 0 26736 0 1 24309
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3265
timestamp 1626908933
transform 1 0 26736 0 1 24309
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1373
timestamp 1626908933
transform 1 0 27024 0 1 24383
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3308
timestamp 1626908933
transform 1 0 27024 0 1 24383
box -29 -23 29 23
use M1M2_PR  M1M2_PR_350
timestamp 1626908933
transform 1 0 27312 0 1 24383
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2317
timestamp 1626908933
transform 1 0 27312 0 1 24383
box -32 -32 32 32
use L1M1_PR  L1M1_PR_372
timestamp 1626908933
transform 1 0 27312 0 1 24383
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2307
timestamp 1626908933
transform 1 0 27312 0 1 24383
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_104
timestamp 1626908933
transform 1 0 27456 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_705
timestamp 1626908933
transform 1 0 27456 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_184
timestamp 1626908933
transform 1 0 27648 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1175
timestamp 1626908933
transform 1 0 27648 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_19
timestamp 1626908933
transform -1 0 27456 0 1 23976
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_7
timestamp 1626908933
transform -1 0 27456 0 1 23976
box -38 -49 1862 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1014
timestamp 1626908933
transform 1 0 28100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_366
timestamp 1626908933
transform 1 0 28100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1014
timestamp 1626908933
transform 1 0 28100 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_366
timestamp 1626908933
transform 1 0 28100 0 1 23976
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_841
timestamp 1626908933
transform 1 0 27744 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_119
timestamp 1626908933
transform 1 0 27744 0 1 23976
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3249
timestamp 1626908933
transform 1 0 29040 0 1 24457
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1282
timestamp 1626908933
transform 1 0 29040 0 1 24457
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1174
timestamp 1626908933
transform 1 0 28896 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_183
timestamp 1626908933
transform 1 0 28896 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_656
timestamp 1626908933
transform 1 0 28512 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_58
timestamp 1626908933
transform 1 0 28512 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_807
timestamp 1626908933
transform 1 0 28992 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_85
timestamp 1626908933
transform 1 0 28992 0 1 23976
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2309
timestamp 1626908933
transform 1 0 29904 0 1 23865
box -32 -32 32 32
use M1M2_PR  M1M2_PR_342
timestamp 1626908933
transform 1 0 29904 0 1 23865
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1160
timestamp 1626908933
transform 1 0 29760 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_704
timestamp 1626908933
transform 1 0 30048 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_559
timestamp 1626908933
transform 1 0 29760 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_103
timestamp 1626908933
transform 1 0 30048 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_448
timestamp 1626908933
transform 1 0 29952 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_91
timestamp 1626908933
transform 1 0 29952 0 1 23976
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2299
timestamp 1626908933
transform 1 0 30192 0 1 23865
box -29 -23 29 23
use L1M1_PR  L1M1_PR_364
timestamp 1626908933
transform 1 0 30192 0 1 23865
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1173
timestamp 1626908933
transform 1 0 30240 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_182
timestamp 1626908933
transform 1 0 30240 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_761
timestamp 1626908933
transform 1 0 30336 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_39
timestamp 1626908933
transform 1 0 30336 0 1 23976
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_990
timestamp 1626908933
transform 1 0 30500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_342
timestamp 1626908933
transform 1 0 30500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_990
timestamp 1626908933
transform 1 0 30500 0 1 23976
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_342
timestamp 1626908933
transform 1 0 30500 0 1 23976
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1172
timestamp 1626908933
transform 1 0 31104 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_181
timestamp 1626908933
transform 1 0 31104 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_727
timestamp 1626908933
transform 1 0 31200 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_5
timestamp 1626908933
transform 1 0 31200 0 1 23976
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3783
timestamp 1626908933
transform 1 0 31920 0 1 23717
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1816
timestamp 1626908933
transform 1 0 31920 0 1 23717
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1923
timestamp 1626908933
transform 1 0 31968 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_932
timestamp 1626908933
transform 1 0 31968 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_102
timestamp 1626908933
transform 1 0 0 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_703
timestamp 1626908933
transform 1 0 0 0 -1 25308
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1543
timestamp 1626908933
transform 1 0 816 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3510
timestamp 1626908933
transform 1 0 816 0 1 24531
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_317
timestamp 1626908933
transform 1 0 500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_965
timestamp 1626908933
transform 1 0 500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_317
timestamp 1626908933
transform 1 0 500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_965
timestamp 1626908933
transform 1 0 500 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_705
timestamp 1626908933
transform 1 0 192 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1427
timestamp 1626908933
transform 1 0 192 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_180
timestamp 1626908933
transform 1 0 960 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1171
timestamp 1626908933
transform 1 0 960 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1126
timestamp 1626908933
transform 1 0 1680 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3093
timestamp 1626908933
transform 1 0 1680 0 1 24753
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1629
timestamp 1626908933
transform 1 0 1584 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3564
timestamp 1626908933
transform 1 0 1584 0 1 24531
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_671
timestamp 1626908933
transform 1 0 1440 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1393
timestamp 1626908933
transform 1 0 1440 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_567
timestamp 1626908933
transform 1 0 1056 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1165
timestamp 1626908933
transform 1 0 1056 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1170
timestamp 1626908933
transform 1 0 2208 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_179
timestamp 1626908933
transform 1 0 2208 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1161
timestamp 1626908933
transform 1 0 2304 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_560
timestamp 1626908933
transform 1 0 2304 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_447
timestamp 1626908933
transform 1 0 2496 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_90
timestamp 1626908933
transform 1 0 2496 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1162
timestamp 1626908933
transform 1 0 2592 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_561
timestamp 1626908933
transform 1 0 2592 0 -1 25308
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_941
timestamp 1626908933
transform 1 0 2900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_293
timestamp 1626908933
transform 1 0 2900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_941
timestamp 1626908933
transform 1 0 2900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_293
timestamp 1626908933
transform 1 0 2900 0 1 24642
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3132
timestamp 1626908933
transform 1 0 2928 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1197
timestamp 1626908933
transform 1 0 2928 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2258
timestamp 1626908933
transform 1 0 3120 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_323
timestamp 1626908933
transform 1 0 3120 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2267
timestamp 1626908933
transform 1 0 3120 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_300
timestamp 1626908933
transform 1 0 3120 0 1 24975
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_178
timestamp 1626908933
transform 1 0 3264 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1169
timestamp 1626908933
transform 1 0 3264 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_123
timestamp 1626908933
transform 1 0 2784 0 -1 25308
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_54
timestamp 1626908933
transform 1 0 2784 0 -1 25308
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_638
timestamp 1626908933
transform 1 0 3360 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1360
timestamp 1626908933
transform 1 0 3360 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_22
timestamp 1626908933
transform -1 0 4704 0 -1 25308
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_9
timestamp 1626908933
transform -1 0 4704 0 -1 25308
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2406
timestamp 1626908933
transform 1 0 4080 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2256
timestamp 1626908933
transform 1 0 4368 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_471
timestamp 1626908933
transform 1 0 4080 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_321
timestamp 1626908933
transform 1 0 4368 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2437
timestamp 1626908933
transform 1 0 4272 0 1 25197
box -32 -32 32 32
use M1M2_PR  M1M2_PR_470
timestamp 1626908933
transform 1 0 4272 0 1 25197
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3214
timestamp 1626908933
transform 1 0 4560 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2167
timestamp 1626908933
transform 1 0 4464 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1279
timestamp 1626908933
transform 1 0 4560 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_232
timestamp 1626908933
transform 1 0 4464 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2394
timestamp 1626908933
transform 1 0 4656 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_459
timestamp 1626908933
transform 1 0 4656 0 1 25049
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2427
timestamp 1626908933
transform 1 0 4656 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_460
timestamp 1626908933
transform 1 0 4656 0 1 25049
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1168
timestamp 1626908933
transform 1 0 4704 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_177
timestamp 1626908933
transform 1 0 4704 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_213
timestamp 1626908933
transform 1 0 4944 0 1 25123
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2180
timestamp 1626908933
transform 1 0 4944 0 1 25123
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_269
timestamp 1626908933
transform 1 0 5300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_917
timestamp 1626908933
transform 1 0 5300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_269
timestamp 1626908933
transform 1 0 5300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_917
timestamp 1626908933
transform 1 0 5300 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_600
timestamp 1626908933
transform 1 0 5184 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1322
timestamp 1626908933
transform 1 0 5184 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_509
timestamp 1626908933
transform 1 0 4800 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1107
timestamp 1626908933
transform 1 0 4800 0 -1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1206
timestamp 1626908933
transform 1 0 5808 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3173
timestamp 1626908933
transform 1 0 5808 0 1 24753
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1281
timestamp 1626908933
transform 1 0 5808 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3216
timestamp 1626908933
transform 1 0 5808 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3209
timestamp 1626908933
transform 1 0 6000 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1274
timestamp 1626908933
transform 1 0 6000 0 1 24753
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3176
timestamp 1626908933
transform 1 0 6000 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1209
timestamp 1626908933
transform 1 0 6000 0 1 24531
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3215
timestamp 1626908933
transform 1 0 6000 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3213
timestamp 1626908933
transform 1 0 6288 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3212
timestamp 1626908933
transform 1 0 6192 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1280
timestamp 1626908933
transform 1 0 6000 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1278
timestamp 1626908933
transform 1 0 6288 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1277
timestamp 1626908933
transform 1 0 6192 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3175
timestamp 1626908933
transform 1 0 6000 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1208
timestamp 1626908933
transform 1 0 6000 0 1 25049
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_702
timestamp 1626908933
transform 1 0 6336 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_101
timestamp 1626908933
transform 1 0 6336 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_58
timestamp 1626908933
transform -1 0 6336 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_120
timestamp 1626908933
transform -1 0 6336 0 -1 25308
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3190
timestamp 1626908933
transform 1 0 6864 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1255
timestamp 1626908933
transform 1 0 6864 0 1 24531
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1294
timestamp 1626908933
transform 1 0 6528 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_572
timestamp 1626908933
transform 1 0 6528 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_89
timestamp 1626908933
transform 1 0 7488 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_446
timestamp 1626908933
transform 1 0 7488 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_100
timestamp 1626908933
transform 1 0 7296 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_701
timestamp 1626908933
transform 1 0 7296 0 -1 25308
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_245
timestamp 1626908933
transform 1 0 7700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_893
timestamp 1626908933
transform 1 0 7700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_245
timestamp 1626908933
transform 1 0 7700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_893
timestamp 1626908933
transform 1 0 7700 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_562
timestamp 1626908933
transform 1 0 7968 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1163
timestamp 1626908933
transform 1 0 7968 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_464
timestamp 1626908933
transform 1 0 7584 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1062
timestamp 1626908933
transform 1 0 7584 0 -1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1193
timestamp 1626908933
transform 1 0 8112 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3160
timestamp 1626908933
transform 1 0 8112 0 1 24531
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1253
timestamp 1626908933
transform 1 0 8208 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3188
timestamp 1626908933
transform 1 0 8208 0 1 24753
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1192
timestamp 1626908933
transform 1 0 8112 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3159
timestamp 1626908933
transform 1 0 8112 0 1 25049
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1254
timestamp 1626908933
transform 1 0 8208 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3189
timestamp 1626908933
transform 1 0 8208 0 1 25049
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_54
timestamp 1626908933
transform -1 0 8544 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_116
timestamp 1626908933
transform -1 0 8544 0 -1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3157
timestamp 1626908933
transform 1 0 8304 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1190
timestamp 1626908933
transform 1 0 8304 0 1 24753
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2390
timestamp 1626908933
transform 1 0 8496 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2156
timestamp 1626908933
transform 1 0 8400 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_455
timestamp 1626908933
transform 1 0 8496 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_221
timestamp 1626908933
transform 1 0 8400 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2420
timestamp 1626908933
transform 1 0 8496 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2169
timestamp 1626908933
transform 1 0 8400 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_453
timestamp 1626908933
transform 1 0 8496 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_202
timestamp 1626908933
transform 1 0 8400 0 1 24975
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_700
timestamp 1626908933
transform 1 0 8544 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_99
timestamp 1626908933
transform 1 0 8544 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_533
timestamp 1626908933
transform 1 0 9120 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1255
timestamp 1626908933
transform 1 0 9120 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_444
timestamp 1626908933
transform 1 0 8736 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1042
timestamp 1626908933
transform 1 0 8736 0 -1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3161
timestamp 1626908933
transform 1 0 9456 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1194
timestamp 1626908933
transform 1 0 9456 0 1 24753
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1167
timestamp 1626908933
transform 1 0 9888 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_176
timestamp 1626908933
transform 1 0 9888 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1015
timestamp 1626908933
transform 1 0 9984 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_417
timestamp 1626908933
transform 1 0 9984 0 -1 25308
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_221
timestamp 1626908933
transform 1 0 10100 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_869
timestamp 1626908933
transform 1 0 10100 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_221
timestamp 1626908933
transform 1 0 10100 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_869
timestamp 1626908933
transform 1 0 10100 0 1 24642
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3211
timestamp 1626908933
transform 1 0 10512 0 1 24901
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2198
timestamp 1626908933
transform 1 0 10608 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1276
timestamp 1626908933
transform 1 0 10512 0 1 24901
box -29 -23 29 23
use L1M1_PR  L1M1_PR_263
timestamp 1626908933
transform 1 0 10608 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2208
timestamp 1626908933
transform 1 0 10608 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_241
timestamp 1626908933
transform 1 0 10608 0 1 24975
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2225
timestamp 1626908933
transform 1 0 10704 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_290
timestamp 1626908933
transform 1 0 10704 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2236
timestamp 1626908933
transform 1 0 10704 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_269
timestamp 1626908933
transform 1 0 10704 0 1 24975
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2423
timestamp 1626908933
transform 1 0 10416 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_488
timestamp 1626908933
transform 1 0 10416 0 1 25049
box -29 -23 29 23
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_10
timestamp 1626908933
transform 1 0 10368 0 -1 25308
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_23
timestamp 1626908933
transform 1 0 10368 0 -1 25308
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2411
timestamp 1626908933
transform 1 0 10992 0 1 24901
box -29 -23 29 23
use L1M1_PR  L1M1_PR_476
timestamp 1626908933
transform 1 0 10992 0 1 24901
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2454
timestamp 1626908933
transform 1 0 10896 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_487
timestamp 1626908933
transform 1 0 10896 0 1 25049
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1166
timestamp 1626908933
transform 1 0 10944 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_175
timestamp 1626908933
transform 1 0 10944 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1214
timestamp 1626908933
transform 1 0 11040 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_492
timestamp 1626908933
transform 1 0 11040 0 -1 25308
box -38 -49 806 715
use M1M2_PR  M1M2_PR_478
timestamp 1626908933
transform 1 0 11472 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1005
timestamp 1626908933
transform 1 0 11088 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2445
timestamp 1626908933
transform 1 0 11472 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2972
timestamp 1626908933
transform 1 0 11088 0 1 24531
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_174
timestamp 1626908933
transform 1 0 11808 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1165
timestamp 1626908933
transform 1 0 11808 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_477
timestamp 1626908933
transform 1 0 11664 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2444
timestamp 1626908933
transform 1 0 11664 0 1 24901
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1069
timestamp 1626908933
transform 1 0 11568 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1256
timestamp 1626908933
transform 1 0 11856 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3004
timestamp 1626908933
transform 1 0 11568 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3191
timestamp 1626908933
transform 1 0 11856 0 1 24753
box -29 -23 29 23
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_4
timestamp 1626908933
transform 1 0 11904 0 -1 25308
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_17
timestamp 1626908933
transform 1 0 11904 0 -1 25308
box -38 -49 614 715
use M1M2_PR  M1M2_PR_2198
timestamp 1626908933
transform 1 0 12048 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_231
timestamp 1626908933
transform 1 0 12048 0 1 24975
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2217
timestamp 1626908933
transform 1 0 12240 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2188
timestamp 1626908933
transform 1 0 12144 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_282
timestamp 1626908933
transform 1 0 12240 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_253
timestamp 1626908933
transform 1 0 12144 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2226
timestamp 1626908933
transform 1 0 12240 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_259
timestamp 1626908933
transform 1 0 12240 0 1 24975
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2418
timestamp 1626908933
transform 1 0 11952 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_483
timestamp 1626908933
transform 1 0 11952 0 1 25049
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_88
timestamp 1626908933
transform 1 0 12480 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_445
timestamp 1626908933
transform 1 0 12480 0 -1 25308
box -38 -49 134 715
use L1M1_PR  L1M1_PR_473
timestamp 1626908933
transform 1 0 12432 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2408
timestamp 1626908933
transform 1 0 12432 0 1 24975
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_197
timestamp 1626908933
transform 1 0 12500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_845
timestamp 1626908933
transform 1 0 12500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_197
timestamp 1626908933
transform 1 0 12500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_845
timestamp 1626908933
transform 1 0 12500 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_358
timestamp 1626908933
transform 1 0 12576 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_956
timestamp 1626908933
transform 1 0 12576 0 -1 25308
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3036
timestamp 1626908933
transform 1 0 13296 0 1 24457
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1101
timestamp 1626908933
transform 1 0 13296 0 1 24457
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1178
timestamp 1626908933
transform 1 0 12960 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_456
timestamp 1626908933
transform 1 0 12960 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_54
timestamp 1626908933
transform 1 0 13728 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_2
timestamp 1626908933
transform 1 0 13728 0 -1 25308
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3040
timestamp 1626908933
transform 1 0 14256 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1105
timestamp 1626908933
transform 1 0 14256 0 1 24531
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3005
timestamp 1626908933
transform 1 0 14448 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1038
timestamp 1626908933
transform 1 0 14448 0 1 24531
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3034
timestamp 1626908933
transform 1 0 14544 0 1 24457
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1099
timestamp 1626908933
transform 1 0 14544 0 1 24457
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3032
timestamp 1626908933
transform 1 0 14064 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1097
timestamp 1626908933
transform 1 0 14064 0 1 24753
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2995
timestamp 1626908933
transform 1 0 14160 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1028
timestamp 1626908933
transform 1 0 14160 0 1 24753
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3035
timestamp 1626908933
transform 1 0 14256 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1100
timestamp 1626908933
transform 1 0 14256 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2999
timestamp 1626908933
transform 1 0 14352 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1032
timestamp 1626908933
transform 1 0 14352 0 1 24901
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3039
timestamp 1626908933
transform 1 0 14448 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1104
timestamp 1626908933
transform 1 0 14448 0 1 25049
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3004
timestamp 1626908933
transform 1 0 14448 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1037
timestamp 1626908933
transform 1 0 14448 0 1 25049
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3601
timestamp 1626908933
transform 1 0 14352 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1666
timestamp 1626908933
transform 1 0 14352 0 1 25197
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_330
timestamp 1626908933
transform 1 0 14496 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_928
timestamp 1626908933
transform 1 0 14496 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_42
timestamp 1626908933
transform 1 0 14112 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_104
timestamp 1626908933
transform 1 0 14112 0 -1 25308
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_821
timestamp 1626908933
transform 1 0 14900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_173
timestamp 1626908933
transform 1 0 14900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_821
timestamp 1626908933
transform 1 0 14900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_173
timestamp 1626908933
transform 1 0 14900 0 1 24642
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3544
timestamp 1626908933
transform 1 0 14928 0 1 25197
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1577
timestamp 1626908933
transform 1 0 14928 0 1 25197
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1142
timestamp 1626908933
transform 1 0 14880 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_420
timestamp 1626908933
transform 1 0 14880 0 -1 25308
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3010
timestamp 1626908933
transform 1 0 15696 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1043
timestamp 1626908933
transform 1 0 15696 0 1 25049
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1164
timestamp 1626908933
transform 1 0 15648 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_173
timestamp 1626908933
transform 1 0 15648 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1111
timestamp 1626908933
transform 1 0 15744 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_389
timestamp 1626908933
transform 1 0 15744 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_110
timestamp 1626908933
transform -1 0 16800 0 -1 25308
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_48
timestamp 1626908933
transform -1 0 16800 0 -1 25308
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3042
timestamp 1626908933
transform 1 0 16560 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1107
timestamp 1626908933
transform 1 0 16560 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3008
timestamp 1626908933
transform 1 0 16464 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1041
timestamp 1626908933
transform 1 0 16464 0 1 24975
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_172
timestamp 1626908933
transform 1 0 16800 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1163
timestamp 1626908933
transform 1 0 16800 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1046
timestamp 1626908933
transform 1 0 16848 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3013
timestamp 1626908933
transform 1 0 16848 0 1 24753
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1110
timestamp 1626908933
transform 1 0 16752 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1115
timestamp 1626908933
transform 1 0 16656 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3045
timestamp 1626908933
transform 1 0 16752 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3050
timestamp 1626908933
transform 1 0 16656 0 1 24753
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_171
timestamp 1626908933
transform 1 0 17280 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_933
timestamp 1626908933
transform 1 0 17376 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1162
timestamp 1626908933
transform 1 0 17280 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1924
timestamp 1626908933
transform 1 0 17376 0 -1 25308
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_149
timestamp 1626908933
transform 1 0 17300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_797
timestamp 1626908933
transform 1 0 17300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_149
timestamp 1626908933
transform 1 0 17300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_797
timestamp 1626908933
transform 1 0 17300 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_286
timestamp 1626908933
transform 1 0 16896 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_884
timestamp 1626908933
transform 1 0 16896 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_87
timestamp 1626908933
transform 1 0 17472 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_444
timestamp 1626908933
transform 1 0 17472 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_170
timestamp 1626908933
transform 1 0 17568 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1161
timestamp 1626908933
transform 1 0 17568 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_169
timestamp 1626908933
transform 1 0 18048 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1160
timestamp 1626908933
transform 1 0 18048 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_350
timestamp 1626908933
transform 1 0 18144 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1072
timestamp 1626908933
transform 1 0 18144 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_263
timestamp 1626908933
transform 1 0 17664 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_861
timestamp 1626908933
transform 1 0 17664 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1159
timestamp 1626908933
transform 1 0 18912 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_168
timestamp 1626908933
transform 1 0 18912 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1045
timestamp 1626908933
transform 1 0 19008 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_323
timestamp 1626908933
transform 1 0 19008 0 -1 25308
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2360
timestamp 1626908933
transform 1 0 19152 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_393
timestamp 1626908933
transform 1 0 19152 0 1 24901
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_773
timestamp 1626908933
transform 1 0 19700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_749
timestamp 1626908933
transform 1 0 22100 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_125
timestamp 1626908933
transform 1 0 19700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_101
timestamp 1626908933
transform 1 0 22100 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_773
timestamp 1626908933
transform 1 0 19700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_749
timestamp 1626908933
transform 1 0 22100 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_125
timestamp 1626908933
transform 1 0 19700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_101
timestamp 1626908933
transform 1 0 22100 0 1 24642
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3399
timestamp 1626908933
transform 1 0 22032 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2298
timestamp 1626908933
transform 1 0 20112 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1464
timestamp 1626908933
transform 1 0 22032 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_363
timestamp 1626908933
transform 1 0 20112 0 1 25197
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3349
timestamp 1626908933
transform 1 0 21648 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2307
timestamp 1626908933
transform 1 0 20208 0 1 25197
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1382
timestamp 1626908933
transform 1 0 21648 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_340
timestamp 1626908933
transform 1 0 20208 0 1 25197
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_65
timestamp 1626908933
transform -1 0 22464 0 -1 25308
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_19
timestamp 1626908933
transform -1 0 22464 0 -1 25308
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3434
timestamp 1626908933
transform 1 0 22416 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1499
timestamp 1626908933
transform 1 0 22416 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3382
timestamp 1626908933
transform 1 0 22512 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1415
timestamp 1626908933
transform 1 0 22512 0 1 24975
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_966
timestamp 1626908933
transform 1 0 22560 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_244
timestamp 1626908933
transform 1 0 22560 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_443
timestamp 1626908933
transform 1 0 22464 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_86
timestamp 1626908933
transform 1 0 22464 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2354
timestamp 1626908933
transform 1 0 23664 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_387
timestamp 1626908933
transform 1 0 23664 0 1 24901
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_699
timestamp 1626908933
transform 1 0 23328 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_98
timestamp 1626908933
transform 1 0 23328 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_753
timestamp 1626908933
transform 1 0 23520 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_155
timestamp 1626908933
transform 1 0 23520 0 -1 25308
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_725
timestamp 1626908933
transform 1 0 24500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_77
timestamp 1626908933
transform 1 0 24500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_725
timestamp 1626908933
transform 1 0 24500 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_77
timestamp 1626908933
transform 1 0 24500 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_936
timestamp 1626908933
transform 1 0 23904 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_214
timestamp 1626908933
transform 1 0 23904 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1158
timestamp 1626908933
transform 1 0 24672 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_167
timestamp 1626908933
transform 1 0 24672 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_728
timestamp 1626908933
transform 1 0 24768 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_130
timestamp 1626908933
transform 1 0 24768 0 -1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3344
timestamp 1626908933
transform 1 0 25488 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1377
timestamp 1626908933
transform 1 0 25488 0 1 25049
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_901
timestamp 1626908933
transform 1 0 25152 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_179
timestamp 1626908933
transform 1 0 25152 0 -1 25308
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3371
timestamp 1626908933
transform 1 0 25776 0 1 24531
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1436
timestamp 1626908933
transform 1 0 25776 0 1 24531
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3320
timestamp 1626908933
transform 1 0 25872 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3319
timestamp 1626908933
transform 1 0 25872 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1353
timestamp 1626908933
transform 1 0 25872 0 1 24531
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1352
timestamp 1626908933
transform 1 0 25872 0 1 24753
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3370
timestamp 1626908933
transform 1 0 26064 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1435
timestamp 1626908933
transform 1 0 26064 0 1 24753
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1925
timestamp 1626908933
transform 1 0 26016 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1157
timestamp 1626908933
transform 1 0 25920 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_934
timestamp 1626908933
transform 1 0 26016 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_166
timestamp 1626908933
transform 1 0 25920 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2304
timestamp 1626908933
transform 1 0 26544 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_337
timestamp 1626908933
transform 1 0 26544 0 1 24975
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3441
timestamp 1626908933
transform 1 0 26352 0 1 25049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1506
timestamp 1626908933
transform 1 0 26352 0 1 25049
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3385
timestamp 1626908933
transform 1 0 26352 0 1 25049
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1418
timestamp 1626908933
transform 1 0 26352 0 1 25049
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3428
timestamp 1626908933
transform 1 0 26448 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1493
timestamp 1626908933
transform 1 0 26448 0 1 25197
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3378
timestamp 1626908933
transform 1 0 26448 0 1 25197
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1411
timestamp 1626908933
transform 1 0 26448 0 1 25197
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_16
timestamp 1626908933
transform 1 0 26112 0 -1 25308
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_41
timestamp 1626908933
transform 1 0 26112 0 -1 25308
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_701
timestamp 1626908933
transform 1 0 26900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_53
timestamp 1626908933
transform 1 0 26900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_701
timestamp 1626908933
transform 1 0 26900 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_53
timestamp 1626908933
transform 1 0 26900 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1156
timestamp 1626908933
transform 1 0 26592 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_165
timestamp 1626908933
transform 1 0 26592 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_862
timestamp 1626908933
transform 1 0 26688 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_140
timestamp 1626908933
transform 1 0 26688 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_698
timestamp 1626908933
transform 1 0 27552 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_97
timestamp 1626908933
transform 1 0 27552 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_442
timestamp 1626908933
transform 1 0 27456 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_85
timestamp 1626908933
transform 1 0 27456 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_2312
timestamp 1626908933
transform 1 0 27792 0 1 25197
box -32 -32 32 32
use M1M2_PR  M1M2_PR_345
timestamp 1626908933
transform 1 0 27792 0 1 25197
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_840
timestamp 1626908933
transform 1 0 27744 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_118
timestamp 1626908933
transform 1 0 27744 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_164
timestamp 1626908933
transform 1 0 28896 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1155
timestamp 1626908933
transform 1 0 28896 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1781
timestamp 1626908933
transform 1 0 28752 0 1 24753
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3748
timestamp 1626908933
transform 1 0 28752 0 1 24753
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_29
timestamp 1626908933
transform 1 0 29300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_677
timestamp 1626908933
transform 1 0 29300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_29
timestamp 1626908933
transform 1 0 29300 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_677
timestamp 1626908933
transform 1 0 29300 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_84
timestamp 1626908933
transform 1 0 28992 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_806
timestamp 1626908933
transform 1 0 28992 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_57
timestamp 1626908933
transform 1 0 28512 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_655
timestamp 1626908933
transform 1 0 28512 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_24
timestamp 1626908933
transform 1 0 30144 0 -1 25308
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_9
timestamp 1626908933
transform 1 0 30144 0 -1 25308
box -38 -49 710 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_625
timestamp 1626908933
transform 1 0 29760 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_27
timestamp 1626908933
transform 1 0 29760 0 -1 25308
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3747
timestamp 1626908933
transform 1 0 30288 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2302
timestamp 1626908933
transform 1 0 30192 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1812
timestamp 1626908933
transform 1 0 30288 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_367
timestamp 1626908933
transform 1 0 30192 0 1 25197
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3793
timestamp 1626908933
transform 1 0 30576 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2340
timestamp 1626908933
transform 1 0 30480 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1858
timestamp 1626908933
transform 1 0 30576 0 1 24975
box -29 -23 29 23
use L1M1_PR  L1M1_PR_405
timestamp 1626908933
transform 1 0 30480 0 1 24975
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3853
timestamp 1626908933
transform 1 0 30576 0 1 24975
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1886
timestamp 1626908933
transform 1 0 30576 0 1 24975
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3728
timestamp 1626908933
transform 1 0 30768 0 1 24753
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1793
timestamp 1626908933
transform 1 0 30768 0 1 24753
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2375
timestamp 1626908933
transform 1 0 30768 0 1 24901
box -32 -32 32 32
use M1M2_PR  M1M2_PR_408
timestamp 1626908933
transform 1 0 30768 0 1 24901
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1154
timestamp 1626908933
transform 1 0 30816 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_163
timestamp 1626908933
transform 1 0 30816 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_24
timestamp 1626908933
transform 1 0 30912 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_746
timestamp 1626908933
transform 1 0 30912 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_84
timestamp 1626908933
transform 1 0 31680 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_441
timestamp 1626908933
transform 1 0 31680 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_563
timestamp 1626908933
transform 1 0 31776 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1164
timestamp 1626908933
transform 1 0 31776 0 -1 25308
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_5
timestamp 1626908933
transform 1 0 31700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_653
timestamp 1626908933
transform 1 0 31700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_5
timestamp 1626908933
transform 1 0 31700 0 1 24642
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_653
timestamp 1626908933
transform 1 0 31700 0 1 24642
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_935
timestamp 1626908933
transform 1 0 31968 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1926
timestamp 1626908933
transform 1 0 31968 0 -1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1817
timestamp 1626908933
transform 1 0 31824 0 1 25123
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3784
timestamp 1626908933
transform 1 0 31824 0 1 25123
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1847
timestamp 1626908933
transform 1 0 48 0 1 25567
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3814
timestamp 1626908933
transform 1 0 48 0 1 25567
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_83
timestamp 1626908933
transform 1 0 288 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_440
timestamp 1626908933
transform 1 0 288 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_936
timestamp 1626908933
transform 1 0 192 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1927
timestamp 1626908933
transform 1 0 192 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_88
timestamp 1626908933
transform 1 0 0 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_564
timestamp 1626908933
transform 1 0 0 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_689
timestamp 1626908933
transform 1 0 0 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1165
timestamp 1626908933
transform 1 0 0 0 1 25308
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_964
timestamp 1626908933
transform 1 0 500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_316
timestamp 1626908933
transform 1 0 500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_964
timestamp 1626908933
transform 1 0 500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_316
timestamp 1626908933
transform 1 0 500 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1188
timestamp 1626908933
transform 1 0 384 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_590
timestamp 1626908933
transform 1 0 384 0 1 25308
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3565
timestamp 1626908933
transform 1 0 816 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1630
timestamp 1626908933
transform 1 0 816 0 1 25641
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3509
timestamp 1626908933
transform 1 0 816 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1542
timestamp 1626908933
transform 1 0 816 0 1 25641
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1146
timestamp 1626908933
transform 1 0 960 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_155
timestamp 1626908933
transform 1 0 960 0 -1 26640
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3664
timestamp 1626908933
transform 1 0 1200 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1729
timestamp 1626908933
transform 1 0 1200 0 1 25641
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1164
timestamp 1626908933
transform 1 0 1056 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_566
timestamp 1626908933
transform 1 0 1056 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_704
timestamp 1626908933
transform 1 0 192 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1426
timestamp 1626908933
transform 1 0 192 0 -1 26640
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_629
timestamp 1626908933
transform 1 0 1700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1277
timestamp 1626908933
transform 1 0 1700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_629
timestamp 1626908933
transform 1 0 1700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1277
timestamp 1626908933
transform 1 0 1700 0 1 25308
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1145
timestamp 1626908933
transform 1 0 2208 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_154
timestamp 1626908933
transform 1 0 2208 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1168
timestamp 1626908933
transform 1 0 2304 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_567
timestamp 1626908933
transform 1 0 2304 0 -1 26640
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3137
timestamp 1626908933
transform 1 0 2448 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1170
timestamp 1626908933
transform 1 0 2448 0 1 25715
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1144
timestamp 1626908933
transform 1 0 2592 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_153
timestamp 1626908933
transform 1 0 2592 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_433
timestamp 1626908933
transform 1 0 2496 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_76
timestamp 1626908933
transform 1 0 2496 0 -1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3610
timestamp 1626908933
transform 1 0 2736 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1643
timestamp 1626908933
transform 1 0 2736 0 1 25641
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_653
timestamp 1626908933
transform 1 0 2688 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_670
timestamp 1626908933
transform 1 0 1440 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1375
timestamp 1626908933
transform 1 0 2688 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1392
timestamp 1626908933
transform 1 0 1440 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_70
timestamp 1626908933
transform 1 0 768 0 1 25308
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_24
timestamp 1626908933
transform 1 0 768 0 1 25308
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_299
timestamp 1626908933
transform 1 0 3120 0 1 25419
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2266
timestamp 1626908933
transform 1 0 3120 0 1 25419
box -32 -32 32 32
use L1M1_PR  L1M1_PR_322
timestamp 1626908933
transform 1 0 3120 0 1 25419
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2257
timestamp 1626908933
transform 1 0 3120 0 1 25419
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_292
timestamp 1626908933
transform 1 0 2900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_940
timestamp 1626908933
transform 1 0 2900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_292
timestamp 1626908933
transform 1 0 2900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_940
timestamp 1626908933
transform 1 0 2900 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_533
timestamp 1626908933
transform 1 0 3456 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_534
timestamp 1626908933
transform 1 0 3456 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1131
timestamp 1626908933
transform 1 0 3456 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1132
timestamp 1626908933
transform 1 0 3456 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_96
timestamp 1626908933
transform 1 0 3840 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_697
timestamp 1626908933
transform 1 0 3840 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_152
timestamp 1626908933
transform 1 0 3840 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_942
timestamp 1626908933
transform 1 0 3936 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1143
timestamp 1626908933
transform 1 0 3840 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1933
timestamp 1626908933
transform 1 0 3936 0 -1 26640
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_605
timestamp 1626908933
transform 1 0 4100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1253
timestamp 1626908933
transform 1 0 4100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_605
timestamp 1626908933
transform 1 0 4100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1253
timestamp 1626908933
transform 1 0 4100 0 1 25308
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_625
timestamp 1626908933
transform 1 0 4032 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1347
timestamp 1626908933
transform 1 0 4032 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_6
timestamp 1626908933
transform -1 0 4608 0 -1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_19
timestamp 1626908933
transform -1 0 4608 0 -1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_95
timestamp 1626908933
transform 1 0 4800 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_696
timestamp 1626908933
transform 1 0 4800 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_82
timestamp 1626908933
transform 1 0 4992 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_439
timestamp 1626908933
transform 1 0 4992 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_94
timestamp 1626908933
transform 1 0 5088 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_695
timestamp 1626908933
transform 1 0 5088 0 1 25308
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_268
timestamp 1626908933
transform 1 0 5300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_916
timestamp 1626908933
transform 1 0 5300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_268
timestamp 1626908933
transform 1 0 5300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_916
timestamp 1626908933
transform 1 0 5300 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_599
timestamp 1626908933
transform 1 0 5280 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_615
timestamp 1626908933
transform 1 0 4608 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1321
timestamp 1626908933
transform 1 0 5280 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1337
timestamp 1626908933
transform 1 0 4608 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_101
timestamp 1626908933
transform 1 0 5376 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_49
timestamp 1626908933
transform 1 0 5376 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_111
timestamp 1626908933
transform 1 0 5760 0 -1 26640
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_42
timestamp 1626908933
transform 1 0 5760 0 -1 26640
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_489
timestamp 1626908933
transform 1 0 6048 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1087
timestamp 1626908933
transform 1 0 6048 0 1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2968
timestamp 1626908933
transform 1 0 6192 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1001
timestamp 1626908933
transform 1 0 6192 0 1 25863
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_688
timestamp 1626908933
transform 1 0 6240 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_87
timestamp 1626908933
transform 1 0 6240 0 -1 26640
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_581
timestamp 1626908933
transform 1 0 6500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1229
timestamp 1626908933
transform 1 0 6500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_581
timestamp 1626908933
transform 1 0 6500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1229
timestamp 1626908933
transform 1 0 6500 0 1 25308
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1072
timestamp 1626908933
transform 1 0 6576 0 1 25419
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3007
timestamp 1626908933
transform 1 0 6576 0 1 25419
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1003
timestamp 1626908933
transform 1 0 6480 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2970
timestamp 1626908933
transform 1 0 6480 0 1 25641
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1067
timestamp 1626908933
transform 1 0 6480 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3002
timestamp 1626908933
transform 1 0 6480 0 1 25641
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_114
timestamp 1626908933
transform 1 0 6432 0 1 25308
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_52
timestamp 1626908933
transform 1 0 6432 0 1 25308
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1081
timestamp 1626908933
transform 1 0 6432 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_483
timestamp 1626908933
transform 1 0 6432 0 -1 26640
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2998
timestamp 1626908933
transform 1 0 6768 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1063
timestamp 1626908933
transform 1 0 6768 0 1 25863
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3177
timestamp 1626908933
transform 1 0 6672 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1210
timestamp 1626908933
transform 1 0 6672 0 1 25715
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1153
timestamp 1626908933
transform 1 0 6720 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_162
timestamp 1626908933
transform 1 0 6720 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1076
timestamp 1626908933
transform 1 0 6816 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_478
timestamp 1626908933
transform 1 0 6816 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_1
timestamp 1626908933
transform 1 0 6816 0 -1 26640
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_9
timestamp 1626908933
transform 1 0 6816 0 -1 26640
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_93
timestamp 1626908933
transform 1 0 7200 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_568
timestamp 1626908933
transform 1 0 7296 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_694
timestamp 1626908933
transform 1 0 7200 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1169
timestamp 1626908933
transform 1 0 7296 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1152
timestamp 1626908933
transform 1 0 7392 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_161
timestamp 1626908933
transform 1 0 7392 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_432
timestamp 1626908933
transform 1 0 7488 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_75
timestamp 1626908933
transform 1 0 7488 0 -1 26640
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_892
timestamp 1626908933
transform 1 0 7700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_244
timestamp 1626908933
transform 1 0 7700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_892
timestamp 1626908933
transform 1 0 7700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_244
timestamp 1626908933
transform 1 0 7700 0 1 25974
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2997
timestamp 1626908933
transform 1 0 7824 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1062
timestamp 1626908933
transform 1 0 7824 0 1 25863
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_99
timestamp 1626908933
transform 1 0 7488 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_47
timestamp 1626908933
transform 1 0 7488 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1061
timestamp 1626908933
transform 1 0 7584 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_463
timestamp 1626908933
transform 1 0 7584 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1934
timestamp 1626908933
transform 1 0 7968 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1928
timestamp 1626908933
transform 1 0 7872 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_943
timestamp 1626908933
transform 1 0 7968 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_937
timestamp 1626908933
transform 1 0 7872 0 1 25308
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3001
timestamp 1626908933
transform 1 0 8112 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1066
timestamp 1626908933
transform 1 0 8112 0 1 25641
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3556
timestamp 1626908933
transform 1 0 8112 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1589
timestamp 1626908933
transform 1 0 8112 0 1 25863
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_101
timestamp 1626908933
transform 1 0 7968 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_39
timestamp 1626908933
transform 1 0 7968 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_85
timestamp 1626908933
transform 1 0 8064 0 -1 26640
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_39
timestamp 1626908933
transform 1 0 8064 0 -1 26640
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_1071
timestamp 1626908933
transform 1 0 8400 0 1 25419
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3006
timestamp 1626908933
transform 1 0 8400 0 1 25419
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_557
timestamp 1626908933
transform 1 0 8900 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1205
timestamp 1626908933
transform 1 0 8900 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_557
timestamp 1626908933
transform 1 0 8900 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1205
timestamp 1626908933
transform 1 0 8900 0 1 25308
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1677
timestamp 1626908933
transform 1 0 8304 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3612
timestamp 1626908933
transform 1 0 8304 0 1 25863
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_119
timestamp 1626908933
transform -1 0 9600 0 1 25308
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_50
timestamp 1626908933
transform -1 0 9600 0 1 25308
box -38 -49 518 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_18
timestamp 1626908933
transform 1 0 8352 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_41
timestamp 1626908933
transform 1 0 8352 0 1 25308
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1089
timestamp 1626908933
transform 1 0 9456 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3056
timestamp 1626908933
transform 1 0 9456 0 1 25863
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1156
timestamp 1626908933
transform 1 0 9456 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3091
timestamp 1626908933
transform 1 0 9456 0 1 25863
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_81
timestamp 1626908933
transform 1 0 9984 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_438
timestamp 1626908933
transform 1 0 9984 0 1 25308
box -38 -49 134 715
use L1M1_PR  L1M1_PR_292
timestamp 1626908933
transform 1 0 9648 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2227
timestamp 1626908933
transform 1 0 9648 0 1 25863
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_48
timestamp 1626908933
transform 1 0 9600 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_100
timestamp 1626908933
transform 1 0 9600 0 1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_271
timestamp 1626908933
transform 1 0 10320 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2238
timestamp 1626908933
transform 1 0 10320 0 1 25863
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_220
timestamp 1626908933
transform 1 0 10100 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_868
timestamp 1626908933
transform 1 0 10100 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_220
timestamp 1626908933
transform 1 0 10100 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_868
timestamp 1626908933
transform 1 0 10100 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_86
timestamp 1626908933
transform 1 0 10752 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_687
timestamp 1626908933
transform 1 0 10752 0 -1 26640
box -38 -49 230 715
use M1M2_PR  M1M2_PR_268
timestamp 1626908933
transform 1 0 10704 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2235
timestamp 1626908933
transform 1 0 10704 0 1 25863
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_19
timestamp 1626908933
transform 1 0 10080 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_42
timestamp 1626908933
transform 1 0 10080 0 1 25308
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2420
timestamp 1626908933
transform 1 0 10896 0 1 25493
box -29 -23 29 23
use L1M1_PR  L1M1_PR_485
timestamp 1626908933
transform 1 0 10896 0 1 25493
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2453
timestamp 1626908933
transform 1 0 10896 0 1 25493
box -32 -32 32 32
use M1M2_PR  M1M2_PR_486
timestamp 1626908933
transform 1 0 10896 0 1 25493
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1929
timestamp 1626908933
transform 1 0 11040 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1142
timestamp 1626908933
transform 1 0 10944 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_938
timestamp 1626908933
transform 1 0 11040 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_151
timestamp 1626908933
transform 1 0 10944 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1166
timestamp 1626908933
transform 1 0 10848 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_565
timestamp 1626908933
transform 1 0 10848 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_491
timestamp 1626908933
transform 1 0 11040 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1213
timestamp 1626908933
transform 1 0 11040 0 -1 26640
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1181
timestamp 1626908933
transform 1 0 11300 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_533
timestamp 1626908933
transform 1 0 11300 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1181
timestamp 1626908933
transform 1 0 11300 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_533
timestamp 1626908933
transform 1 0 11300 0 1 25308
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2971
timestamp 1626908933
transform 1 0 11088 0 1 25419
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1004
timestamp 1626908933
transform 1 0 11088 0 1 25419
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1282
timestamp 1626908933
transform 1 0 11280 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3217
timestamp 1626908933
transform 1 0 11280 0 1 25715
box -29 -23 29 23
use M1M2_PR  M1M2_PR_263
timestamp 1626908933
transform 1 0 11472 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2230
timestamp 1626908933
transform 1 0 11472 0 1 25641
box -32 -32 32 32
use L1M1_PR  L1M1_PR_256
timestamp 1626908933
transform 1 0 11376 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_285
timestamp 1626908933
transform 1 0 11472 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2191
timestamp 1626908933
transform 1 0 11376 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2220
timestamp 1626908933
transform 1 0 11472 0 1 25641
box -29 -23 29 23
use M1M2_PR  M1M2_PR_476
timestamp 1626908933
transform 1 0 11664 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2443
timestamp 1626908933
transform 1 0 11664 0 1 25641
box -32 -32 32 32
use L1M1_PR  L1M1_PR_475
timestamp 1626908933
transform 1 0 11664 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2410
timestamp 1626908933
transform 1 0 11664 0 1 25641
box -29 -23 29 23
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_25
timestamp 1626908933
transform 1 0 11136 0 1 25308
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_12
timestamp 1626908933
transform 1 0 11136 0 1 25308
box -38 -49 614 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_983
timestamp 1626908933
transform 1 0 11712 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_385
timestamp 1626908933
transform 1 0 11712 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1141
timestamp 1626908933
transform 1 0 12000 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_150
timestamp 1626908933
transform 1 0 12000 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_686
timestamp 1626908933
transform 1 0 11808 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_85
timestamp 1626908933
transform 1 0 11808 0 -1 26640
box -38 -49 230 715
use L1M1_PR  L1M1_PR_2190
timestamp 1626908933
transform 1 0 12240 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_255
timestamp 1626908933
transform 1 0 12240 0 1 25715
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1167
timestamp 1626908933
transform 1 0 12096 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_566
timestamp 1626908933
transform 1 0 12096 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_974
timestamp 1626908933
transform 1 0 12096 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_376
timestamp 1626908933
transform 1 0 12096 0 -1 26640
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_196
timestamp 1626908933
transform 1 0 12500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_844
timestamp 1626908933
transform 1 0 12500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_196
timestamp 1626908933
transform 1 0 12500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_844
timestamp 1626908933
transform 1 0 12500 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_74
timestamp 1626908933
transform 1 0 12480 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_431
timestamp 1626908933
transform 1 0 12480 0 -1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_233
timestamp 1626908933
transform 1 0 13008 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2200
timestamp 1626908933
transform 1 0 13008 0 1 25715
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_42
timestamp 1626908933
transform 1 0 13344 0 -1 26640
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_103
timestamp 1626908933
transform 1 0 13344 0 -1 26640
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1720
timestamp 1626908933
transform 1 0 13488 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3687
timestamp 1626908933
transform 1 0 13488 0 1 25715
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_509
timestamp 1626908933
transform 1 0 13700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1157
timestamp 1626908933
transform 1 0 13700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_509
timestamp 1626908933
transform 1 0 13700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1157
timestamp 1626908933
transform 1 0 13700 0 1 25308
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_437
timestamp 1626908933
transform 1 0 13632 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_455
timestamp 1626908933
transform 1 0 12576 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1159
timestamp 1626908933
transform 1 0 13632 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1177
timestamp 1626908933
transform 1 0 12576 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_86
timestamp 1626908933
transform -1 0 14976 0 1 25308
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_40
timestamp 1626908933
transform -1 0 14976 0 1 25308
box -38 -49 2726 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_149
timestamp 1626908933
transform 1 0 14400 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1140
timestamp 1626908933
transform 1 0 14400 0 -1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1036
timestamp 1626908933
transform 1 0 14448 0 1 25419
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1613
timestamp 1626908933
transform 1 0 14544 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3003
timestamp 1626908933
transform 1 0 14448 0 1 25419
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3580
timestamp 1626908933
transform 1 0 14544 0 1 25641
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1705
timestamp 1626908933
transform 1 0 14544 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3640
timestamp 1626908933
transform 1 0 14544 0 1 25641
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_329
timestamp 1626908933
transform 1 0 14496 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_927
timestamp 1626908933
transform 1 0 14496 0 -1 26640
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_820
timestamp 1626908933
transform 1 0 14900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_172
timestamp 1626908933
transform 1 0 14900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_820
timestamp 1626908933
transform 1 0 14900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_172
timestamp 1626908933
transform 1 0 14900 0 1 25974
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2202
timestamp 1626908933
transform 1 0 14832 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_235
timestamp 1626908933
transform 1 0 14832 0 1 25715
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3600
timestamp 1626908933
transform 1 0 14928 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1665
timestamp 1626908933
transform 1 0 14928 0 1 25641
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3543
timestamp 1626908933
transform 1 0 14928 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1576
timestamp 1626908933
transform 1 0 14928 0 1 25641
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_437
timestamp 1626908933
transform 1 0 14976 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_80
timestamp 1626908933
transform 1 0 14976 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_160
timestamp 1626908933
transform 1 0 15456 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1151
timestamp 1626908933
transform 1 0 15456 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_419
timestamp 1626908933
transform 1 0 14880 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1141
timestamp 1626908933
transform 1 0 14880 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_315
timestamp 1626908933
transform 1 0 15072 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_913
timestamp 1626908933
transform 1 0 15072 0 1 25308
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1133
timestamp 1626908933
transform 1 0 16100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_485
timestamp 1626908933
transform 1 0 16100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1133
timestamp 1626908933
transform 1 0 16100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_485
timestamp 1626908933
transform 1 0 16100 0 1 25308
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3037
timestamp 1626908933
transform 1 0 16272 0 1 25419
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1102
timestamp 1626908933
transform 1 0 16272 0 1 25419
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3002
timestamp 1626908933
transform 1 0 16176 0 1 25419
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1035
timestamp 1626908933
transform 1 0 16176 0 1 25419
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_106
timestamp 1626908933
transform 1 0 16320 0 1 25308
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_45
timestamp 1626908933
transform 1 0 16320 0 1 25308
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_403
timestamp 1626908933
transform 1 0 15552 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1125
timestamp 1626908933
transform 1 0 15552 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_303
timestamp 1626908933
transform 1 0 15648 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_901
timestamp 1626908933
transform 1 0 15648 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_29
timestamp 1626908933
transform -1 0 16608 0 -1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_68
timestamp 1626908933
transform -1 0 16608 0 -1 26640
box -38 -49 614 715
use L1M1_PR  L1M1_PR_3043
timestamp 1626908933
transform 1 0 16464 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1108
timestamp 1626908933
transform 1 0 16464 0 1 25863
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3007
timestamp 1626908933
transform 1 0 16464 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1040
timestamp 1626908933
transform 1 0 16464 0 1 25863
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_92
timestamp 1626908933
transform 1 0 16608 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_693
timestamp 1626908933
transform 1 0 16608 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_148
timestamp 1626908933
transform 1 0 16608 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1139
timestamp 1626908933
transform 1 0 16608 0 -1 26640
box -38 -49 134 715
use L1M1_PR  L1M1_PR_257
timestamp 1626908933
transform 1 0 16656 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2192
timestamp 1626908933
transform 1 0 16656 0 1 25715
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_148
timestamp 1626908933
transform 1 0 17300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_796
timestamp 1626908933
transform 1 0 17300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_148
timestamp 1626908933
transform 1 0 17300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_796
timestamp 1626908933
transform 1 0 17300 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_376
timestamp 1626908933
transform 1 0 16704 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_377
timestamp 1626908933
transform 1 0 16800 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1098
timestamp 1626908933
transform 1 0 16704 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1099
timestamp 1626908933
transform 1 0 16800 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_73
timestamp 1626908933
transform 1 0 17472 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_430
timestamp 1626908933
transform 1 0 17472 0 -1 26640
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1824
timestamp 1626908933
transform 1 0 18000 0 1 25567
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3759
timestamp 1626908933
transform 1 0 18000 0 1 25567
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_261
timestamp 1626908933
transform 1 0 17568 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_262
timestamp 1626908933
transform 1 0 17568 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_859
timestamp 1626908933
transform 1 0 17568 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_860
timestamp 1626908933
transform 1 0 17568 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_1
timestamp 1626908933
transform 1 0 17952 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_53
timestamp 1626908933
transform 1 0 17952 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_2
timestamp 1626908933
transform 1 0 17952 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_8
timestamp 1626908933
transform 1 0 17952 0 1 25308
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_461
timestamp 1626908933
transform 1 0 18500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1109
timestamp 1626908933
transform 1 0 18500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_461
timestamp 1626908933
transform 1 0 18500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1109
timestamp 1626908933
transform 1 0 18500 0 1 25308
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1306
timestamp 1626908933
transform 1 0 18960 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1311
timestamp 1626908933
transform 1 0 18480 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3273
timestamp 1626908933
transform 1 0 18960 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3278
timestamp 1626908933
transform 1 0 18480 0 1 25641
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1381
timestamp 1626908933
transform 1 0 18672 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1391
timestamp 1626908933
transform 1 0 18480 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3316
timestamp 1626908933
transform 1 0 18672 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3326
timestamp 1626908933
transform 1 0 18480 0 1 25641
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_335
timestamp 1626908933
transform 1 0 18720 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1057
timestamp 1626908933
transform 1 0 18720 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_50
timestamp 1626908933
transform 1 0 18336 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_102
timestamp 1626908933
transform 1 0 18336 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_1
timestamp 1626908933
transform 1 0 18720 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_7
timestamp 1626908933
transform 1 0 18720 0 -1 26640
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_772
timestamp 1626908933
transform 1 0 19700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_124
timestamp 1626908933
transform 1 0 19700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_772
timestamp 1626908933
transform 1 0 19700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_124
timestamp 1626908933
transform 1 0 19700 0 1 25974
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3259
timestamp 1626908933
transform 1 0 19440 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1292
timestamp 1626908933
transform 1 0 19440 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3257
timestamp 1626908933
transform 1 0 19920 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1290
timestamp 1626908933
transform 1 0 19920 0 1 25863
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1930
timestamp 1626908933
transform 1 0 19872 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_939
timestamp 1626908933
transform 1 0 19872 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_685
timestamp 1626908933
transform 1 0 19872 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_84
timestamp 1626908933
transform 1 0 19872 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_436
timestamp 1626908933
transform 1 0 19968 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_79
timestamp 1626908933
transform 1 0 19968 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_825
timestamp 1626908933
transform 1 0 19488 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_824
timestamp 1626908933
transform 1 0 19488 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_227
timestamp 1626908933
transform 1 0 19488 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_226
timestamp 1626908933
transform 1 0 19488 0 -1 26640
box -38 -49 422 715
use M1M2_PR  M1M2_PR_339
timestamp 1626908933
transform 1 0 20208 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1285
timestamp 1626908933
transform 1 0 20400 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2306
timestamp 1626908933
transform 1 0 20208 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3252
timestamp 1626908933
transform 1 0 20400 0 1 25715
box -32 -32 32 32
use L1M1_PR  L1M1_PR_362
timestamp 1626908933
transform 1 0 20208 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1378
timestamp 1626908933
transform 1 0 20496 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2297
timestamp 1626908933
transform 1 0 20208 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3313
timestamp 1626908933
transform 1 0 20496 0 1 25715
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_305
timestamp 1626908933
transform 1 0 20064 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1027
timestamp 1626908933
transform 1 0 20064 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_201
timestamp 1626908933
transform 1 0 20928 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_799
timestamp 1626908933
transform 1 0 20928 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_147
timestamp 1626908933
transform 1 0 20832 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1138
timestamp 1626908933
transform 1 0 20832 0 -1 26640
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_437
timestamp 1626908933
transform 1 0 20900 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1085
timestamp 1626908933
transform 1 0 20900 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_437
timestamp 1626908933
transform 1 0 20900 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1085
timestamp 1626908933
transform 1 0 20900 0 1 25308
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3376
timestamp 1626908933
transform 1 0 21744 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3312
timestamp 1626908933
transform 1 0 21552 0 1 25715
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1441
timestamp 1626908933
transform 1 0 21744 0 1 25863
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1377
timestamp 1626908933
transform 1 0 21552 0 1 25715
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3326
timestamp 1626908933
transform 1 0 21648 0 1 25863
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1359
timestamp 1626908933
transform 1 0 21648 0 1 25863
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_748
timestamp 1626908933
transform 1 0 22100 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_100
timestamp 1626908933
transform 1 0 22100 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_748
timestamp 1626908933
transform 1 0 22100 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_100
timestamp 1626908933
transform 1 0 22100 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1150
timestamp 1626908933
transform 1 0 21888 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_159
timestamp 1626908933
transform 1 0 21888 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_780
timestamp 1626908933
transform 1 0 22080 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_182
timestamp 1626908933
transform 1 0 22080 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_267
timestamp 1626908933
transform 1 0 21984 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_280
timestamp 1626908933
transform 1 0 21312 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_989
timestamp 1626908933
transform 1 0 21984 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1002
timestamp 1626908933
transform 1 0 21312 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_22
timestamp 1626908933
transform 1 0 20064 0 1 25308
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_10
timestamp 1626908933
transform 1 0 20064 0 1 25308
box -38 -49 1862 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_72
timestamp 1626908933
transform 1 0 22464 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_429
timestamp 1626908933
transform 1 0 22464 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_569
timestamp 1626908933
transform 1 0 22560 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1170
timestamp 1626908933
transform 1 0 22560 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_158
timestamp 1626908933
transform 1 0 22752 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1149
timestamp 1626908933
transform 1 0 22752 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_169
timestamp 1626908933
transform 1 0 22848 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_767
timestamp 1626908933
transform 1 0 22848 0 1 25308
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1284
timestamp 1626908933
transform 1 0 23184 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3251
timestamp 1626908933
transform 1 0 23184 0 1 25715
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_413
timestamp 1626908933
transform 1 0 23300 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1061
timestamp 1626908933
transform 1 0 23300 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_413
timestamp 1626908933
transform 1 0 23300 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1061
timestamp 1626908933
transform 1 0 23300 0 1 25308
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_230
timestamp 1626908933
transform 1 0 23232 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_952
timestamp 1626908933
transform 1 0 23232 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_91
timestamp 1626908933
transform 1 0 24000 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_692
timestamp 1626908933
transform 1 0 24000 0 1 25308
box -38 -49 230 715
use M1M2_PR  M1M2_PR_386
timestamp 1626908933
transform 1 0 23664 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2353
timestamp 1626908933
transform 1 0 23664 0 1 25715
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_129
timestamp 1626908933
transform 1 0 24768 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_727
timestamp 1626908933
transform 1 0 24768 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_83
timestamp 1626908933
transform 1 0 24576 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_684
timestamp 1626908933
transform 1 0 24576 0 -1 26640
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_76
timestamp 1626908933
transform 1 0 24500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_724
timestamp 1626908933
transform 1 0 24500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_76
timestamp 1626908933
transform 1 0 24500 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_724
timestamp 1626908933
transform 1 0 24500 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_199
timestamp 1626908933
transform 1 0 24192 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_921
timestamp 1626908933
transform 1 0 24192 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_21
timestamp 1626908933
transform 1 0 22752 0 -1 26640
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_9
timestamp 1626908933
transform 1 0 22752 0 -1 26640
box -38 -49 1862 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_78
timestamp 1626908933
transform 1 0 24960 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_435
timestamp 1626908933
transform 1 0 24960 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_940
timestamp 1626908933
transform 1 0 25056 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1931
timestamp 1626908933
transform 1 0 25056 0 1 25308
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1376
timestamp 1626908933
transform 1 0 25488 0 1 25641
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3343
timestamp 1626908933
transform 1 0 25488 0 1 25641
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1494
timestamp 1626908933
transform 1 0 25200 0 1 25567
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3429
timestamp 1626908933
transform 1 0 25200 0 1 25567
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1037
timestamp 1626908933
transform 1 0 25700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_389
timestamp 1626908933
transform 1 0 25700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1037
timestamp 1626908933
transform 1 0 25700 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_389
timestamp 1626908933
transform 1 0 25700 0 1 25308
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3392
timestamp 1626908933
transform 1 0 25584 0 1 25641
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1457
timestamp 1626908933
transform 1 0 25584 0 1 25641
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_683
timestamp 1626908933
transform 1 0 25920 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_82
timestamp 1626908933
transform 1 0 25920 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_700
timestamp 1626908933
transform 1 0 26112 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_102
timestamp 1626908933
transform 1 0 26112 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_178
timestamp 1626908933
transform 1 0 25152 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_900
timestamp 1626908933
transform 1 0 25152 0 -1 26640
box -38 -49 806 715
use M1M2_PR  M1M2_PR_380
timestamp 1626908933
transform 1 0 26544 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1410
timestamp 1626908933
transform 1 0 26448 0 1 25567
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2347
timestamp 1626908933
transform 1 0 26544 0 1 25715
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3377
timestamp 1626908933
transform 1 0 26448 0 1 25567
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_52
timestamp 1626908933
transform 1 0 26900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_700
timestamp 1626908933
transform 1 0 26900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_52
timestamp 1626908933
transform 1 0 26900 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_700
timestamp 1626908933
transform 1 0 26900 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_71
timestamp 1626908933
transform 1 0 27456 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_428
timestamp 1626908933
transform 1 0 27456 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_570
timestamp 1626908933
transform 1 0 27264 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1171
timestamp 1626908933
transform 1 0 27264 0 -1 26640
box -38 -49 230 715
use M1M2_PR  M1M2_PR_349
timestamp 1626908933
transform 1 0 27312 0 1 25419
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2316
timestamp 1626908933
transform 1 0 27312 0 1 25419
box -32 -32 32 32
use L1M1_PR  L1M1_PR_371
timestamp 1626908933
transform 1 0 27504 0 1 25419
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2306
timestamp 1626908933
transform 1 0 27504 0 1 25419
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_150
timestamp 1626908933
transform 1 0 26496 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_872
timestamp 1626908933
transform 1 0 26496 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_20
timestamp 1626908933
transform 1 0 27552 0 -1 26640
box -38 -49 1862 715
use sky130_fd_sc_hs__fa_2  sky130_fd_sc_hs__fa_2_8
timestamp 1626908933
transform 1 0 27552 0 -1 26640
box -38 -49 1862 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_47
timestamp 1626908933
transform 1 0 25152 0 1 25308
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_1
timestamp 1626908933
transform 1 0 25152 0 1 25308
box -38 -49 2726 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_90
timestamp 1626908933
transform 1 0 27840 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_691
timestamp 1626908933
transform 1 0 27840 0 1 25308
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_365
timestamp 1626908933
transform 1 0 28100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1013
timestamp 1626908933
transform 1 0 28100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_365
timestamp 1626908933
transform 1 0 28100 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1013
timestamp 1626908933
transform 1 0 28100 0 1 25308
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_106
timestamp 1626908933
transform 1 0 28416 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_828
timestamp 1626908933
transform 1 0 28416 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_73
timestamp 1626908933
transform 1 0 28032 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_671
timestamp 1626908933
transform 1 0 28032 0 1 25308
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_676
timestamp 1626908933
transform 1 0 29300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_28
timestamp 1626908933
transform 1 0 29300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_676
timestamp 1626908933
transform 1 0 29300 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_28
timestamp 1626908933
transform 1 0 29300 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_793
timestamp 1626908933
transform 1 0 29184 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_71
timestamp 1626908933
transform 1 0 29184 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_81
timestamp 1626908933
transform 1 0 29376 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_682
timestamp 1626908933
transform 1 0 29376 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_146
timestamp 1626908933
transform 1 0 29568 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1137
timestamp 1626908933
transform 1 0 29568 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_77
timestamp 1626908933
transform 1 0 29952 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_434
timestamp 1626908933
transform 1 0 29952 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_89
timestamp 1626908933
transform 1 0 30048 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_690
timestamp 1626908933
transform 1 0 30048 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_70
timestamp 1626908933
transform 1 0 29664 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_792
timestamp 1626908933
transform 1 0 29664 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1148
timestamp 1626908933
transform 1 0 30240 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_157
timestamp 1626908933
transform 1 0 30240 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_760
timestamp 1626908933
transform 1 0 30336 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_38
timestamp 1626908933
transform 1 0 30336 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_145
timestamp 1626908933
transform 1 0 30432 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1136
timestamp 1626908933
transform 1 0 30432 0 -1 26640
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_341
timestamp 1626908933
transform 1 0 30500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_989
timestamp 1626908933
transform 1 0 30500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_341
timestamp 1626908933
transform 1 0 30500 0 1 25308
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_989
timestamp 1626908933
transform 1 0 30500 0 1 25308
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_156
timestamp 1626908933
transform 1 0 31104 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1147
timestamp 1626908933
transform 1 0 31104 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_4
timestamp 1626908933
transform 1 0 31200 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_23
timestamp 1626908933
transform 1 0 30912 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_726
timestamp 1626908933
transform 1 0 31200 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_745
timestamp 1626908933
transform 1 0 30912 0 -1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_19
timestamp 1626908933
transform 1 0 30528 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_617
timestamp 1626908933
transform 1 0 30528 0 -1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_70
timestamp 1626908933
transform 1 0 31680 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_427
timestamp 1626908933
transform 1 0 31680 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_571
timestamp 1626908933
transform 1 0 31776 0 -1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1172
timestamp 1626908933
transform 1 0 31776 0 -1 26640
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_4
timestamp 1626908933
transform 1 0 31700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_652
timestamp 1626908933
transform 1 0 31700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_4
timestamp 1626908933
transform 1 0 31700 0 1 25974
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_652
timestamp 1626908933
transform 1 0 31700 0 1 25974
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_941
timestamp 1626908933
transform 1 0 31968 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_944
timestamp 1626908933
transform 1 0 31968 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1932
timestamp 1626908933
transform 1 0 31968 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1935
timestamp 1626908933
transform 1 0 31968 0 -1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_69
timestamp 1626908933
transform 1 0 288 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_426
timestamp 1626908933
transform 1 0 288 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_572
timestamp 1626908933
transform 1 0 0 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1173
timestamp 1626908933
transform 1 0 0 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_945
timestamp 1626908933
transform 1 0 192 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1936
timestamp 1626908933
transform 1 0 192 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1846
timestamp 1626908933
transform 1 0 48 0 1 26455
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3813
timestamp 1626908933
transform 1 0 48 0 1 26455
box -32 -32 32 32
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_37
timestamp 1626908933
transform 1 0 1152 0 1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_76
timestamp 1626908933
transform 1 0 1152 0 1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_692
timestamp 1626908933
transform 1 0 384 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1414
timestamp 1626908933
transform 1 0 384 0 1 26640
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1276
timestamp 1626908933
transform 1 0 1700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_628
timestamp 1626908933
transform 1 0 1700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1276
timestamp 1626908933
transform 1 0 1700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_628
timestamp 1626908933
transform 1 0 1700 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_681
timestamp 1626908933
transform 1 0 1728 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_80
timestamp 1626908933
transform 1 0 1728 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1151
timestamp 1626908933
transform 1 0 1920 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_553
timestamp 1626908933
transform 1 0 1920 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_67
timestamp 1626908933
transform 1 0 2304 0 1 26640
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_21
timestamp 1626908933
transform 1 0 2304 0 1 26640
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_472
timestamp 1626908933
transform 1 0 3984 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2407
timestamp 1626908933
transform 1 0 3984 0 1 26085
box -29 -23 29 23
use M1M2_PR  M1M2_PR_296
timestamp 1626908933
transform 1 0 3888 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2263
timestamp 1626908933
transform 1 0 3888 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_298
timestamp 1626908933
transform 1 0 3504 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2265
timestamp 1626908933
transform 1 0 3504 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_295
timestamp 1626908933
transform 1 0 3888 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2262
timestamp 1626908933
transform 1 0 3888 0 1 26751
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_604
timestamp 1626908933
transform 1 0 4100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1252
timestamp 1626908933
transform 1 0 4100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_604
timestamp 1626908933
transform 1 0 4100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1252
timestamp 1626908933
transform 1 0 4100 0 1 26640
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2436
timestamp 1626908933
transform 1 0 4272 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_469
timestamp 1626908933
transform 1 0 4272 0 1 26085
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2253
timestamp 1626908933
transform 1 0 4272 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_318
timestamp 1626908933
transform 1 0 4272 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3200
timestamp 1626908933
transform 1 0 4464 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2163
timestamp 1626908933
transform 1 0 4368 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1265
timestamp 1626908933
transform 1 0 4464 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_228
timestamp 1626908933
transform 1 0 4368 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2395
timestamp 1626908933
transform 1 0 4560 0 1 26381
box -29 -23 29 23
use L1M1_PR  L1M1_PR_460
timestamp 1626908933
transform 1 0 4560 0 1 26381
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_68
timestamp 1626908933
transform 1 0 4992 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_425
timestamp 1626908933
transform 1 0 4992 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_211
timestamp 1626908933
transform 1 0 5040 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_212
timestamp 1626908933
transform 1 0 4944 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_459
timestamp 1626908933
transform 1 0 4656 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2178
timestamp 1626908933
transform 1 0 5040 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2179
timestamp 1626908933
transform 1 0 4944 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2426
timestamp 1626908933
transform 1 0 4656 0 1 26381
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_500
timestamp 1626908933
transform 1 0 5088 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1098
timestamp 1626908933
transform 1 0 5088 0 1 26640
box -38 -49 422 715
use M1M2_PR  M1M2_PR_210
timestamp 1626908933
transform 1 0 5520 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2177
timestamp 1626908933
transform 1 0 5520 0 1 26233
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_82
timestamp 1626908933
transform -1 0 8160 0 1 26640
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_36
timestamp 1626908933
transform -1 0 8160 0 1 26640
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_2165
timestamp 1626908933
transform 1 0 5712 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_230
timestamp 1626908933
transform 1 0 5712 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3003
timestamp 1626908933
transform 1 0 6096 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1068
timestamp 1626908933
transform 1 0 6096 0 1 26085
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2482
timestamp 1626908933
transform 1 0 6288 0 1 26159
box -32 -32 32 32
use M1M2_PR  M1M2_PR_515
timestamp 1626908933
transform 1 0 6288 0 1 26159
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1228
timestamp 1626908933
transform 1 0 6500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_580
timestamp 1626908933
transform 1 0 6500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1228
timestamp 1626908933
transform 1 0 6500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_580
timestamp 1626908933
transform 1 0 6500 0 1 26640
box -100 -49 100 49
use M1M2_PR  M1M2_PR_2969
timestamp 1626908933
transform 1 0 6480 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1002
timestamp 1626908933
transform 1 0 6480 0 1 26085
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3199
timestamp 1626908933
transform 1 0 6960 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2445
timestamp 1626908933
transform 1 0 6960 0 1 26159
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1264
timestamp 1626908933
transform 1 0 6960 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_510
timestamp 1626908933
transform 1 0 6960 0 1 26159
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3198
timestamp 1626908933
transform 1 0 7152 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1263
timestamp 1626908933
transform 1 0 7152 0 1 26307
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3712
timestamp 1626908933
transform 1 0 7824 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3168
timestamp 1626908933
transform 1 0 7920 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1745
timestamp 1626908933
transform 1 0 7824 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1201
timestamp 1626908933
transform 1 0 7920 0 1 26307
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3581
timestamp 1626908933
transform 1 0 8112 0 1 26381
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1646
timestamp 1626908933
transform 1 0 8112 0 1 26381
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_680
timestamp 1626908933
transform 1 0 8160 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_79
timestamp 1626908933
transform 1 0 8160 0 1 26640
box -38 -49 230 715
use M1M2_PR  M1M2_PR_3524
timestamp 1626908933
transform 1 0 8304 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3523
timestamp 1626908933
transform 1 0 8304 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1557
timestamp 1626908933
transform 1 0 8304 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1556
timestamp 1626908933
transform 1 0 8304 0 1 26751
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1135
timestamp 1626908933
transform 1 0 8352 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_144
timestamp 1626908933
transform 1 0 8352 0 1 26640
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3650
timestamp 1626908933
transform 1 0 8496 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1715
timestamp 1626908933
transform 1 0 8496 0 1 26307
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3594
timestamp 1626908933
transform 1 0 8688 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1627
timestamp 1626908933
transform 1 0 8688 0 1 26307
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_556
timestamp 1626908933
transform 1 0 8900 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1204
timestamp 1626908933
transform 1 0 8900 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_556
timestamp 1626908933
transform 1 0 8900 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1204
timestamp 1626908933
transform 1 0 8900 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_546
timestamp 1626908933
transform 1 0 8448 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1268
timestamp 1626908933
transform 1 0 8448 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_109
timestamp 1626908933
transform -1 0 9600 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_47
timestamp 1626908933
transform -1 0 9600 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_103
timestamp 1626908933
transform 1 0 9600 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_51
timestamp 1626908933
transform 1 0 9600 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_424
timestamp 1626908933
transform 1 0 9984 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_67
timestamp 1626908933
transform 1 0 9984 0 1 26640
box -38 -49 134 715
use L1M1_PR  L1M1_PR_2226
timestamp 1626908933
transform 1 0 10320 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_291
timestamp 1626908933
transform 1 0 10320 0 1 26085
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2237
timestamp 1626908933
transform 1 0 10320 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_270
timestamp 1626908933
transform 1 0 10320 0 1 26085
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1014
timestamp 1626908933
transform 1 0 10080 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_416
timestamp 1626908933
transform 1 0 10080 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1229
timestamp 1626908933
transform 1 0 10464 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_507
timestamp 1626908933
transform 1 0 10464 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_573
timestamp 1626908933
transform 1 0 11232 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1174
timestamp 1626908933
transform 1 0 11232 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_946
timestamp 1626908933
transform 1 0 11424 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1937
timestamp 1626908933
transform 1 0 11424 0 1 26640
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_532
timestamp 1626908933
transform 1 0 11300 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1180
timestamp 1626908933
transform 1 0 11300 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_532
timestamp 1626908933
transform 1 0 11300 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1180
timestamp 1626908933
transform 1 0 11300 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_7
timestamp 1626908933
transform 1 0 11520 0 1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_20
timestamp 1626908933
transform 1 0 11520 0 1 26640
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_78
timestamp 1626908933
transform 1 0 12096 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_679
timestamp 1626908933
transform 1 0 12096 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_143
timestamp 1626908933
transform 1 0 12288 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1134
timestamp 1626908933
transform 1 0 12288 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_258
timestamp 1626908933
transform 1 0 12240 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2225
timestamp 1626908933
transform 1 0 12240 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_255
timestamp 1626908933
transform 1 0 12720 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2222
timestamp 1626908933
transform 1 0 12720 0 1 26233
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_468
timestamp 1626908933
transform 1 0 12384 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1190
timestamp 1626908933
transform 1 0 12384 0 1 26640
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3036
timestamp 1626908933
transform 1 0 13296 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1069
timestamp 1626908933
transform 1 0 13296 0 1 26381
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3071
timestamp 1626908933
transform 1 0 13392 0 1 26381
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1136
timestamp 1626908933
transform 1 0 13392 0 1 26381
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3077
timestamp 1626908933
transform 1 0 13584 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2214
timestamp 1626908933
transform 1 0 13584 0 1 26381
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1142
timestamp 1626908933
transform 1 0 13584 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_279
timestamp 1626908933
transform 1 0 13584 0 1 26381
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1133
timestamp 1626908933
transform 1 0 13536 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_142
timestamp 1626908933
transform 1 0 13536 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_351
timestamp 1626908933
transform 1 0 13152 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_949
timestamp 1626908933
transform 1 0 13152 0 1 26640
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1156
timestamp 1626908933
transform 1 0 13700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_508
timestamp 1626908933
transform 1 0 13700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1156
timestamp 1626908933
transform 1 0 13700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_508
timestamp 1626908933
transform 1 0 13700 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1158
timestamp 1626908933
transform 1 0 13632 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_436
timestamp 1626908933
transform 1 0 13632 0 1 26640
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3043
timestamp 1626908933
transform 1 0 13872 0 1 26529
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1076
timestamp 1626908933
transform 1 0 13872 0 1 26529
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_678
timestamp 1626908933
transform 1 0 14400 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_77
timestamp 1626908933
transform 1 0 14400 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_926
timestamp 1626908933
transform 1 0 14592 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_328
timestamp 1626908933
transform 1 0 14592 0 1 26640
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2205
timestamp 1626908933
transform 1 0 14736 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_238
timestamp 1626908933
transform 1 0 14736 0 1 26307
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1132
timestamp 1626908933
transform 1 0 15456 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_141
timestamp 1626908933
transform 1 0 15456 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_912
timestamp 1626908933
transform 1 0 15072 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_314
timestamp 1626908933
transform 1 0 15072 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_423
timestamp 1626908933
transform 1 0 14976 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_66
timestamp 1626908933
transform 1 0 14976 0 1 26640
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1132
timestamp 1626908933
transform 1 0 16100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_484
timestamp 1626908933
transform 1 0 16100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1132
timestamp 1626908933
transform 1 0 16100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_484
timestamp 1626908933
transform 1 0 16100 0 1 26640
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2193
timestamp 1626908933
transform 1 0 16080 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_258
timestamp 1626908933
transform 1 0 16080 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3038
timestamp 1626908933
transform 1 0 16176 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1103
timestamp 1626908933
transform 1 0 16176 0 1 26085
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3001
timestamp 1626908933
transform 1 0 16176 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1034
timestamp 1626908933
transform 1 0 16176 0 1 26085
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1131
timestamp 1626908933
transform 1 0 16320 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_140
timestamp 1626908933
transform 1 0 16320 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_402
timestamp 1626908933
transform 1 0 15552 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1124
timestamp 1626908933
transform 1 0 15552 0 1 26640
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3599
timestamp 1626908933
transform 1 0 16560 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3044
timestamp 1626908933
transform 1 0 16368 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1664
timestamp 1626908933
transform 1 0 16560 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1109
timestamp 1626908933
transform 1 0 16368 0 1 26307
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3006
timestamp 1626908933
transform 1 0 16464 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1039
timestamp 1626908933
transform 1 0 16464 0 1 26307
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_892
timestamp 1626908933
transform 1 0 16416 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_294
timestamp 1626908933
transform 1 0 16416 0 1 26640
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3542
timestamp 1626908933
transform 1 0 16752 0 1 26529
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1575
timestamp 1626908933
transform 1 0 16752 0 1 26529
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1097
timestamp 1626908933
transform 1 0 16800 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_375
timestamp 1626908933
transform 1 0 16800 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1130
timestamp 1626908933
transform 1 0 17568 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1129
timestamp 1626908933
transform 1 0 18048 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_139
timestamp 1626908933
transform 1 0 17568 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_138
timestamp 1626908933
transform 1 0 18048 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_858
timestamp 1626908933
transform 1 0 17664 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_260
timestamp 1626908933
transform 1 0 17664 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1071
timestamp 1626908933
transform 1 0 18144 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_349
timestamp 1626908933
transform 1 0 18144 0 1 26640
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1310
timestamp 1626908933
transform 1 0 18480 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3277
timestamp 1626908933
transform 1 0 18480 0 1 26307
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_460
timestamp 1626908933
transform 1 0 18500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1108
timestamp 1626908933
transform 1 0 18500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_460
timestamp 1626908933
transform 1 0 18500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1108
timestamp 1626908933
transform 1 0 18500 0 1 26640
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1823
timestamp 1626908933
transform 1 0 18576 0 1 26455
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3758
timestamp 1626908933
transform 1 0 18576 0 1 26455
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_76
timestamp 1626908933
transform 1 0 18912 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_677
timestamp 1626908933
transform 1 0 18912 0 1 26640
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1389
timestamp 1626908933
transform 1 0 19056 0 1 26307
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3324
timestamp 1626908933
transform 1 0 19056 0 1 26307
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_137
timestamp 1626908933
transform 1 0 19104 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1128
timestamp 1626908933
transform 1 0 19104 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1044
timestamp 1626908933
transform 1 0 19200 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_322
timestamp 1626908933
transform 1 0 19200 0 1 26640
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1291
timestamp 1626908933
transform 1 0 19440 0 1 26085
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3258
timestamp 1626908933
transform 1 0 19440 0 1 26085
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1382
timestamp 1626908933
transform 1 0 19440 0 1 26085
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3317
timestamp 1626908933
transform 1 0 19440 0 1 26085
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_65
timestamp 1626908933
transform 1 0 19968 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_422
timestamp 1626908933
transform 1 0 19968 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_75
timestamp 1626908933
transform 1 0 20064 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_676
timestamp 1626908933
transform 1 0 20064 0 1 26640
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1289
timestamp 1626908933
transform 1 0 19920 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3256
timestamp 1626908933
transform 1 0 19920 0 1 26307
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_947
timestamp 1626908933
transform 1 0 20640 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1938
timestamp 1626908933
transform 1 0 20640 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1305
timestamp 1626908933
transform 1 0 20688 0 1 26529
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3272
timestamp 1626908933
transform 1 0 20688 0 1 26529
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_436
timestamp 1626908933
transform 1 0 20900 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1084
timestamp 1626908933
transform 1 0 20900 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_436
timestamp 1626908933
transform 1 0 20900 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1084
timestamp 1626908933
transform 1 0 20900 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_214
timestamp 1626908933
transform 1 0 20256 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_812
timestamp 1626908933
transform 1 0 20256 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_13
timestamp 1626908933
transform -1 0 21216 0 1 26640
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_38
timestamp 1626908933
transform -1 0 21216 0 1 26640
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1127
timestamp 1626908933
transform 1 0 21216 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_136
timestamp 1626908933
transform 1 0 21216 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1001
timestamp 1626908933
transform 1 0 21312 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_279
timestamp 1626908933
transform 1 0 21312 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_779
timestamp 1626908933
transform 1 0 22080 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_181
timestamp 1626908933
transform 1 0 22080 0 1 26640
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2301
timestamp 1626908933
transform 1 0 22896 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_366
timestamp 1626908933
transform 1 0 22896 0 1 26233
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3381
timestamp 1626908933
transform 1 0 22512 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1414
timestamp 1626908933
transform 1 0 22512 0 1 26751
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1126
timestamp 1626908933
transform 1 0 22464 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_135
timestamp 1626908933
transform 1 0 22464 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_965
timestamp 1626908933
transform 1 0 22560 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_243
timestamp 1626908933
transform 1 0 22560 0 1 26640
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3311
timestamp 1626908933
transform 1 0 23184 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1376
timestamp 1626908933
transform 1 0 23184 0 1 26233
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3250
timestamp 1626908933
transform 1 0 23184 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1283
timestamp 1626908933
transform 1 0 23184 0 1 26233
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1060
timestamp 1626908933
transform 1 0 23300 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_412
timestamp 1626908933
transform 1 0 23300 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1060
timestamp 1626908933
transform 1 0 23300 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_412
timestamp 1626908933
transform 1 0 23300 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_675
timestamp 1626908933
transform 1 0 23328 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_74
timestamp 1626908933
transform 1 0 23328 0 1 26640
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1357
timestamp 1626908933
transform 1 0 23760 0 1 26529
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3324
timestamp 1626908933
transform 1 0 23760 0 1 26529
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_154
timestamp 1626908933
transform 1 0 23520 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_752
timestamp 1626908933
transform 1 0 23520 0 1 26640
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3374
timestamp 1626908933
transform 1 0 24432 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3310
timestamp 1626908933
transform 1 0 24240 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1439
timestamp 1626908933
transform 1 0 24432 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1375
timestamp 1626908933
transform 1 0 24240 0 1 26233
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2311
timestamp 1626908933
transform 1 0 23952 0 1 26159
box -32 -32 32 32
use M1M2_PR  M1M2_PR_344
timestamp 1626908933
transform 1 0 23952 0 1 26159
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_935
timestamp 1626908933
transform 1 0 23904 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_213
timestamp 1626908933
transform 1 0 23904 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1939
timestamp 1626908933
transform 1 0 24864 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_948
timestamp 1626908933
transform 1 0 24864 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1175
timestamp 1626908933
transform 1 0 24672 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_574
timestamp 1626908933
transform 1 0 24672 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_64
timestamp 1626908933
transform 1 0 24960 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_421
timestamp 1626908933
transform 1 0 24960 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_134
timestamp 1626908933
transform 1 0 25056 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1125
timestamp 1626908933
transform 1 0 25056 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1287
timestamp 1626908933
transform 1 0 25200 0 1 26307
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3254
timestamp 1626908933
transform 1 0 25200 0 1 26307
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_388
timestamp 1626908933
transform 1 0 25700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1036
timestamp 1626908933
transform 1 0 25700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_388
timestamp 1626908933
transform 1 0 25700 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1036
timestamp 1626908933
transform 1 0 25700 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_177
timestamp 1626908933
transform 1 0 25152 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_899
timestamp 1626908933
transform 1 0 25152 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_674
timestamp 1626908933
transform 1 0 25920 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_73
timestamp 1626908933
transform 1 0 25920 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_699
timestamp 1626908933
transform 1 0 26112 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_101
timestamp 1626908933
transform 1 0 26112 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_871
timestamp 1626908933
transform 1 0 26496 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_149
timestamp 1626908933
transform 1 0 26496 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1124
timestamp 1626908933
transform 1 0 27264 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_133
timestamp 1626908933
transform 1 0 27264 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_679
timestamp 1626908933
transform 1 0 27360 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_81
timestamp 1626908933
transform 1 0 27360 0 1 26640
box -38 -49 422 715
use M1M2_PR  M1M2_PR_347
timestamp 1626908933
transform 1 0 27696 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2314
timestamp 1626908933
transform 1 0 27696 0 1 26233
box -32 -32 32 32
use L1M1_PR  L1M1_PR_368
timestamp 1626908933
transform 1 0 27696 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1374
timestamp 1626908933
transform 1 0 27984 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2303
timestamp 1626908933
transform 1 0 27696 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3309
timestamp 1626908933
transform 1 0 27984 0 1 26233
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_364
timestamp 1626908933
transform 1 0 28100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1012
timestamp 1626908933
transform 1 0 28100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_364
timestamp 1626908933
transform 1 0 28100 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1012
timestamp 1626908933
transform 1 0 28100 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_117
timestamp 1626908933
transform 1 0 27744 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_839
timestamp 1626908933
transform 1 0 27744 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_132
timestamp 1626908933
transform 1 0 28896 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1123
timestamp 1626908933
transform 1 0 28896 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1819
timestamp 1626908933
transform 1 0 28560 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3786
timestamp 1626908933
transform 1 0 28560 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1281
timestamp 1626908933
transform 1 0 29040 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1355
timestamp 1626908933
transform 1 0 29136 0 1 26529
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3248
timestamp 1626908933
transform 1 0 29040 0 1 26233
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3322
timestamp 1626908933
transform 1 0 29136 0 1 26529
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1372
timestamp 1626908933
transform 1 0 29040 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1437
timestamp 1626908933
transform 1 0 29232 0 1 26529
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3307
timestamp 1626908933
transform 1 0 29040 0 1 26233
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3372
timestamp 1626908933
transform 1 0 29232 0 1 26529
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_83
timestamp 1626908933
transform 1 0 28992 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_805
timestamp 1626908933
transform 1 0 28992 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_56
timestamp 1626908933
transform 1 0 28512 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_654
timestamp 1626908933
transform 1 0 28512 0 1 26640
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1940
timestamp 1626908933
transform 1 0 29856 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1122
timestamp 1626908933
transform 1 0 29760 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_949
timestamp 1626908933
transform 1 0 29856 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_131
timestamp 1626908933
transform 1 0 29760 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_673
timestamp 1626908933
transform 1 0 30048 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_72
timestamp 1626908933
transform 1 0 30048 0 1 26640
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_420
timestamp 1626908933
transform 1 0 29952 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_63
timestamp 1626908933
transform 1 0 29952 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1121
timestamp 1626908933
transform 1 0 30240 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_130
timestamp 1626908933
transform 1 0 30240 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_759
timestamp 1626908933
transform 1 0 30336 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_37
timestamp 1626908933
transform 1 0 30336 0 1 26640
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_340
timestamp 1626908933
transform 1 0 30500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_988
timestamp 1626908933
transform 1 0 30500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_340
timestamp 1626908933
transform 1 0 30500 0 1 26640
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_988
timestamp 1626908933
transform 1 0 30500 0 1 26640
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_129
timestamp 1626908933
transform 1 0 31104 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1120
timestamp 1626908933
transform 1 0 31104 0 1 26640
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1822
timestamp 1626908933
transform 1 0 31248 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3789
timestamp 1626908933
transform 1 0 31248 0 1 26751
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_3
timestamp 1626908933
transform 1 0 31200 0 1 26640
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_725
timestamp 1626908933
transform 1 0 31200 0 1 26640
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3788
timestamp 1626908933
transform 1 0 32016 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3785
timestamp 1626908933
transform 1 0 31920 0 1 26381
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1821
timestamp 1626908933
transform 1 0 32016 0 1 26751
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1818
timestamp 1626908933
transform 1 0 31920 0 1 26381
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1941
timestamp 1626908933
transform 1 0 31968 0 1 26640
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_950
timestamp 1626908933
transform 1 0 31968 0 1 26640
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_963
timestamp 1626908933
transform 1 0 500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_315
timestamp 1626908933
transform 1 0 500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_963
timestamp 1626908933
transform 1 0 500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_315
timestamp 1626908933
transform 1 0 500 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_672
timestamp 1626908933
transform 1 0 0 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_71
timestamp 1626908933
transform 1 0 0 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1425
timestamp 1626908933
transform 1 0 192 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_703
timestamp 1626908933
transform 1 0 192 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_128
timestamp 1626908933
transform 1 0 960 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1119
timestamp 1626908933
transform 1 0 960 0 -1 27972
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1632
timestamp 1626908933
transform 1 0 1200 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3567
timestamp 1626908933
transform 1 0 1200 0 1 26899
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1123
timestamp 1626908933
transform 1 0 1296 0 1 26973
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3090
timestamp 1626908933
transform 1 0 1296 0 1 26973
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1192
timestamp 1626908933
transform 1 0 1584 0 1 27195
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1195
timestamp 1626908933
transform 1 0 1392 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3127
timestamp 1626908933
transform 1 0 1584 0 1 27195
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3130
timestamp 1626908933
transform 1 0 1392 0 1 26973
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_669
timestamp 1626908933
transform 1 0 1440 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1391
timestamp 1626908933
transform 1 0 1440 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_565
timestamp 1626908933
transform 1 0 1056 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1163
timestamp 1626908933
transform 1 0 1056 0 -1 27972
box -38 -49 422 715
use L1M1_PR  L1M1_PR_320
timestamp 1626908933
transform 1 0 1776 0 1 26751
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2255
timestamp 1626908933
transform 1 0 1776 0 1 26751
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_127
timestamp 1626908933
transform 1 0 2208 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1118
timestamp 1626908933
transform 1 0 2208 0 -1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1120
timestamp 1626908933
transform 1 0 1968 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1121
timestamp 1626908933
transform 1 0 1968 0 1 27195
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3087
timestamp 1626908933
transform 1 0 1968 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3088
timestamp 1626908933
transform 1 0 1968 0 1 27195
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_62
timestamp 1626908933
transform 1 0 2496 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_419
timestamp 1626908933
transform 1 0 2496 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_575
timestamp 1626908933
transform 1 0 2304 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1176
timestamp 1626908933
transform 1 0 2304 0 -1 27972
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1169
timestamp 1626908933
transform 1 0 2448 0 1 27047
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3136
timestamp 1626908933
transform 1 0 2448 0 1 27047
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1631
timestamp 1626908933
transform 1 0 2352 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3566
timestamp 1626908933
transform 1 0 2352 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3663
timestamp 1626908933
transform 1 0 2736 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1728
timestamp 1626908933
transform 1 0 2736 0 1 26973
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3609
timestamp 1626908933
transform 1 0 2736 0 1 26825
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1642
timestamp 1626908933
transform 1 0 2736 0 1 26825
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1177
timestamp 1626908933
transform 1 0 2592 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_576
timestamp 1626908933
transform 1 0 2592 0 -1 27972
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_939
timestamp 1626908933
transform 1 0 2900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_291
timestamp 1626908933
transform 1 0 2900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_939
timestamp 1626908933
transform 1 0 2900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_291
timestamp 1626908933
transform 1 0 2900 0 1 27306
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3125
timestamp 1626908933
transform 1 0 2832 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1190
timestamp 1626908933
transform 1 0 2832 0 1 27417
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1942
timestamp 1626908933
transform 1 0 2784 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_951
timestamp 1626908933
transform 1 0 2784 0 -1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3135
timestamp 1626908933
transform 1 0 3120 0 1 27047
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1168
timestamp 1626908933
transform 1 0 3120 0 1 27047
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_671
timestamp 1626908933
transform 1 0 3168 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_70
timestamp 1626908933
transform 1 0 3168 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_98
timestamp 1626908933
transform 1 0 2880 0 -1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_37
timestamp 1626908933
transform 1 0 2880 0 -1 27972
box -38 -49 326 715
use M1M2_PR  M1M2_PR_297
timestamp 1626908933
transform 1 0 3504 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2264
timestamp 1626908933
transform 1 0 3504 0 1 27417
box -32 -32 32 32
use L1M1_PR  L1M1_PR_319
timestamp 1626908933
transform 1 0 3216 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2254
timestamp 1626908933
transform 1 0 3216 0 1 27417
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_637
timestamp 1626908933
transform 1 0 3360 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1359
timestamp 1626908933
transform 1 0 3360 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_24
timestamp 1626908933
transform 1 0 4320 0 -1 27972
box -38 -49 614 715
use sky130_fd_sc_hs__a22oi_1  sky130_fd_sc_hs__a22oi_1_11
timestamp 1626908933
transform 1 0 4320 0 -1 27972
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2396
timestamp 1626908933
transform 1 0 4176 0 1 27491
box -29 -23 29 23
use L1M1_PR  L1M1_PR_461
timestamp 1626908933
transform 1 0 4176 0 1 27491
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2435
timestamp 1626908933
transform 1 0 4272 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_468
timestamp 1626908933
transform 1 0 4272 0 1 27417
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_670
timestamp 1626908933
transform 1 0 4128 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_69
timestamp 1626908933
transform 1 0 4128 0 -1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_317
timestamp 1626908933
transform 1 0 4656 0 1 26751
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2252
timestamp 1626908933
transform 1 0 4656 0 1 26751
box -29 -23 29 23
use M1M2_PR  M1M2_PR_458
timestamp 1626908933
transform 1 0 4656 0 1 27491
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2425
timestamp 1626908933
transform 1 0 4656 0 1 27491
box -32 -32 32 32
use L1M1_PR  L1M1_PR_467
timestamp 1626908933
transform 1 0 4944 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2402
timestamp 1626908933
transform 1 0 4944 0 1 27417
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_267
timestamp 1626908933
transform 1 0 5300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_915
timestamp 1626908933
transform 1 0 5300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_267
timestamp 1626908933
transform 1 0 5300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_915
timestamp 1626908933
transform 1 0 5300 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_598
timestamp 1626908933
transform 1 0 5280 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1320
timestamp 1626908933
transform 1 0 5280 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_0
timestamp 1626908933
transform 1 0 4896 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_52
timestamp 1626908933
transform 1 0 4896 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_577
timestamp 1626908933
transform 1 0 6048 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1178
timestamp 1626908933
transform 1 0 6048 0 -1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_231
timestamp 1626908933
transform 1 0 5616 0 1 26751
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2166
timestamp 1626908933
transform 1 0 5616 0 1 26751
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_49
timestamp 1626908933
transform -1 0 6528 0 -1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_110
timestamp 1626908933
transform -1 0 6528 0 -1 27972
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1164
timestamp 1626908933
transform 1 0 6384 0 1 27195
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3131
timestamp 1626908933
transform 1 0 6384 0 1 27195
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_20
timestamp 1626908933
transform 1 0 6528 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_43
timestamp 1626908933
transform 1 0 6528 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_578
timestamp 1626908933
transform 1 0 7296 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1179
timestamp 1626908933
transform 1 0 7296 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_61
timestamp 1626908933
transform 1 0 7488 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_418
timestamp 1626908933
transform 1 0 7488 0 -1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1632
timestamp 1626908933
transform 1 0 7536 0 1 26973
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3599
timestamp 1626908933
transform 1 0 7536 0 1 26973
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_243
timestamp 1626908933
transform 1 0 7700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_891
timestamp 1626908933
transform 1 0 7700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_243
timestamp 1626908933
transform 1 0 7700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_891
timestamp 1626908933
transform 1 0 7700 0 1 27306
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1744
timestamp 1626908933
transform 1 0 7824 0 1 27047
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3711
timestamp 1626908933
transform 1 0 7824 0 1 27047
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1719
timestamp 1626908933
transform 1 0 7728 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3654
timestamp 1626908933
transform 1 0 7728 0 1 26973
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1200
timestamp 1626908933
transform 1 0 8016 0 1 27047
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1588
timestamp 1626908933
transform 1 0 8112 0 1 26973
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3167
timestamp 1626908933
transform 1 0 8016 0 1 27047
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3555
timestamp 1626908933
transform 1 0 8112 0 1 26973
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1678
timestamp 1626908933
transform 1 0 8112 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3613
timestamp 1626908933
transform 1 0 8112 0 1 26973
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_56
timestamp 1626908933
transform 1 0 7584 0 -1 27972
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_10
timestamp 1626908933
transform 1 0 7584 0 -1 27972
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_3597
timestamp 1626908933
transform 1 0 8304 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3593
timestamp 1626908933
transform 1 0 8688 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1630
timestamp 1626908933
transform 1 0 8304 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1626
timestamp 1626908933
transform 1 0 8688 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1094
timestamp 1626908933
transform 1 0 9264 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3061
timestamp 1626908933
transform 1 0 9264 0 1 26899
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1159
timestamp 1626908933
transform 1 0 9264 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3094
timestamp 1626908933
transform 1 0 9264 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1645
timestamp 1626908933
transform 1 0 9360 0 1 26751
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3580
timestamp 1626908933
transform 1 0 9360 0 1 26751
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1090
timestamp 1626908933
transform 1 0 9840 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3057
timestamp 1626908933
transform 1 0 9840 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1088
timestamp 1626908933
transform 1 0 9456 0 1 26973
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3055
timestamp 1626908933
transform 1 0 9456 0 1 26973
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1155
timestamp 1626908933
transform 1 0 9456 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3090
timestamp 1626908933
transform 1 0 9456 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1153
timestamp 1626908933
transform 1 0 9648 0 1 27195
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3088
timestamp 1626908933
transform 1 0 9648 0 1 27195
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1086
timestamp 1626908933
transform 1 0 9840 0 1 27195
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3053
timestamp 1626908933
transform 1 0 9840 0 1 27195
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1085
timestamp 1626908933
transform 1 0 9840 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3052
timestamp 1626908933
transform 1 0 9840 0 1 27417
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_867
timestamp 1626908933
transform 1 0 10100 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_219
timestamp 1626908933
transform 1 0 10100 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_867
timestamp 1626908933
transform 1 0 10100 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_219
timestamp 1626908933
transform 1 0 10100 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1117
timestamp 1626908933
transform 1 0 10272 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_126
timestamp 1626908933
transform 1 0 10272 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1228
timestamp 1626908933
transform 1 0 10368 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_506
timestamp 1626908933
transform 1 0 10368 0 -1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2452
timestamp 1626908933
transform 1 0 10896 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_485
timestamp 1626908933
transform 1 0 10896 0 1 26899
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_41
timestamp 1626908933
transform 1 0 11136 0 -1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_102
timestamp 1626908933
transform 1 0 11136 0 -1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_68
timestamp 1626908933
transform 1 0 11424 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_669
timestamp 1626908933
transform 1 0 11424 0 -1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_289
timestamp 1626908933
transform 1 0 11472 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1151
timestamp 1626908933
transform 1 0 11280 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2224
timestamp 1626908933
transform 1 0 11472 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3086
timestamp 1626908933
transform 1 0 11280 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2419
timestamp 1626908933
transform 1 0 11568 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_484
timestamp 1626908933
transform 1 0 11568 0 1 26899
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1116
timestamp 1626908933
transform 1 0 11616 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_125
timestamp 1626908933
transform 1 0 11616 0 -1 27972
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3197
timestamp 1626908933
transform 1 0 11664 0 1 27047
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2195
timestamp 1626908933
transform 1 0 11760 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1262
timestamp 1626908933
transform 1 0 11664 0 1 27047
box -29 -23 29 23
use L1M1_PR  L1M1_PR_260
timestamp 1626908933
transform 1 0 11760 0 1 26973
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2442
timestamp 1626908933
transform 1 0 11664 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_475
timestamp 1626908933
transform 1 0 11664 0 1 26899
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2223
timestamp 1626908933
transform 1 0 11856 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_288
timestamp 1626908933
transform 1 0 11856 0 1 26973
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2234
timestamp 1626908933
transform 1 0 11856 0 1 26973
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2233
timestamp 1626908933
transform 1 0 11856 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_267
timestamp 1626908933
transform 1 0 11856 0 1 26973
box -32 -32 32 32
use M1M2_PR  M1M2_PR_266
timestamp 1626908933
transform 1 0 11856 0 1 27417
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_478
timestamp 1626908933
transform 1 0 11712 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1200
timestamp 1626908933
transform 1 0 11712 0 -1 27972
box -38 -49 806 715
use L1M1_PR  L1M1_PR_474
timestamp 1626908933
transform 1 0 12048 0 1 26973
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2409
timestamp 1626908933
transform 1 0 12048 0 1 26973
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_195
timestamp 1626908933
transform 1 0 12500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_843
timestamp 1626908933
transform 1 0 12500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_195
timestamp 1626908933
transform 1 0 12500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_843
timestamp 1626908933
transform 1 0 12500 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_60
timestamp 1626908933
transform 1 0 12480 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_417
timestamp 1626908933
transform 1 0 12480 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_67
timestamp 1626908933
transform 1 0 12576 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_668
timestamp 1626908933
transform 1 0 12576 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_71
timestamp 1626908933
transform -1 0 14112 0 -1 27972
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_32
timestamp 1626908933
transform -1 0 14112 0 -1 27972
box -38 -49 614 715
use M1M2_PR  M1M2_PR_3035
timestamp 1626908933
transform 1 0 13296 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1068
timestamp 1626908933
transform 1 0 13296 0 1 27417
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1176
timestamp 1626908933
transform 1 0 12768 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_454
timestamp 1626908933
transform 1 0 12768 0 -1 27972
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3070
timestamp 1626908933
transform 1 0 13680 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1135
timestamp 1626908933
transform 1 0 13680 0 1 27417
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_66
timestamp 1626908933
transform 1 0 14112 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_667
timestamp 1626908933
transform 1 0 14112 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_340
timestamp 1626908933
transform 1 0 14304 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_938
timestamp 1626908933
transform 1 0 14304 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_952
timestamp 1626908933
transform 1 0 14688 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1943
timestamp 1626908933
transform 1 0 14688 0 -1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_236
timestamp 1626908933
transform 1 0 14736 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_237
timestamp 1626908933
transform 1 0 14736 0 1 27047
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2203
timestamp 1626908933
transform 1 0 14736 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2204
timestamp 1626908933
transform 1 0 14736 0 1 27047
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_171
timestamp 1626908933
transform 1 0 14900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_819
timestamp 1626908933
transform 1 0 14900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_171
timestamp 1626908933
transform 1 0 14900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_819
timestamp 1626908933
transform 1 0 14900 0 1 27306
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2194
timestamp 1626908933
transform 1 0 15216 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_259
timestamp 1626908933
transform 1 0 15216 0 1 27417
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_78
timestamp 1626908933
transform -1 0 17472 0 -1 27972
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_32
timestamp 1626908933
transform -1 0 17472 0 -1 27972
box -38 -49 2726 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_795
timestamp 1626908933
transform 1 0 17300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_147
timestamp 1626908933
transform 1 0 17300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_795
timestamp 1626908933
transform 1 0 17300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_147
timestamp 1626908933
transform 1 0 17300 0 1 27306
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3541
timestamp 1626908933
transform 1 0 16752 0 1 27491
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1574
timestamp 1626908933
transform 1 0 16752 0 1 27491
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_59
timestamp 1626908933
transform 1 0 17472 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_416
timestamp 1626908933
transform 1 0 17472 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_124
timestamp 1626908933
transform 1 0 17568 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1115
timestamp 1626908933
transform 1 0 17568 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_123
timestamp 1626908933
transform 1 0 18048 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1114
timestamp 1626908933
transform 1 0 18048 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_348
timestamp 1626908933
transform 1 0 18144 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1070
timestamp 1626908933
transform 1 0 18144 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_259
timestamp 1626908933
transform 1 0 17664 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_857
timestamp 1626908933
transform 1 0 17664 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1113
timestamp 1626908933
transform 1 0 18912 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_122
timestamp 1626908933
transform 1 0 18912 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_834
timestamp 1626908933
transform 1 0 19008 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_236
timestamp 1626908933
transform 1 0 19008 0 -1 27972
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_771
timestamp 1626908933
transform 1 0 19700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_123
timestamp 1626908933
transform 1 0 19700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_771
timestamp 1626908933
transform 1 0 19700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_123
timestamp 1626908933
transform 1 0 19700 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1112
timestamp 1626908933
transform 1 0 20160 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_121
timestamp 1626908933
transform 1 0 20160 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1043
timestamp 1626908933
transform 1 0 19392 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_321
timestamp 1626908933
transform 1 0 19392 0 -1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1431
timestamp 1626908933
transform 1 0 20976 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3398
timestamp 1626908933
transform 1 0 20976 0 1 26899
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1500
timestamp 1626908933
transform 1 0 20880 0 1 26751
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1516
timestamp 1626908933
transform 1 0 20976 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3435
timestamp 1626908933
transform 1 0 20880 0 1 26751
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3451
timestamp 1626908933
transform 1 0 20976 0 1 26899
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_295
timestamp 1626908933
transform 1 0 20640 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1017
timestamp 1626908933
transform 1 0 20640 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_213
timestamp 1626908933
transform 1 0 20256 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_811
timestamp 1626908933
transform 1 0 20256 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_65
timestamp 1626908933
transform 1 0 21408 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_666
timestamp 1626908933
transform 1 0 21408 0 -1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1442
timestamp 1626908933
transform 1 0 21168 0 1 26899
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3377
timestamp 1626908933
transform 1 0 21168 0 1 26899
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_120
timestamp 1626908933
transform 1 0 21600 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1111
timestamp 1626908933
transform 1 0 21600 0 -1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1358
timestamp 1626908933
transform 1 0 21648 0 1 26899
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3325
timestamp 1626908933
transform 1 0 21648 0 1 26899
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_266
timestamp 1626908933
transform 1 0 21696 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_988
timestamp 1626908933
transform 1 0 21696 0 -1 27972
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_747
timestamp 1626908933
transform 1 0 22100 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_99
timestamp 1626908933
transform 1 0 22100 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_747
timestamp 1626908933
transform 1 0 22100 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_99
timestamp 1626908933
transform 1 0 22100 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_58
timestamp 1626908933
transform 1 0 22464 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_415
timestamp 1626908933
transform 1 0 22464 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_64
timestamp 1626908933
transform 1 0 22560 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_665
timestamp 1626908933
transform 1 0 22560 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_168
timestamp 1626908933
transform 1 0 22848 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_766
timestamp 1626908933
transform 1 0 22848 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_119
timestamp 1626908933
transform 1 0 22752 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1110
timestamp 1626908933
transform 1 0 22752 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_10
timestamp 1626908933
transform -1 0 23712 0 -1 27972
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_35
timestamp 1626908933
transform -1 0 23712 0 -1 27972
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_63
timestamp 1626908933
transform 1 0 23712 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_664
timestamp 1626908933
transform 1 0 23712 0 -1 27972
box -38 -49 230 715
use M1M2_PR  M1M2_PR_343
timestamp 1626908933
transform 1 0 23952 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1356
timestamp 1626908933
transform 1 0 23760 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2310
timestamp 1626908933
transform 1 0 23952 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3323
timestamp 1626908933
transform 1 0 23760 0 1 27417
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1440
timestamp 1626908933
transform 1 0 23760 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3375
timestamp 1626908933
transform 1 0 23760 0 1 27417
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_75
timestamp 1626908933
transform 1 0 24500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_723
timestamp 1626908933
transform 1 0 24500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_75
timestamp 1626908933
transform 1 0 24500 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_723
timestamp 1626908933
transform 1 0 24500 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_212
timestamp 1626908933
transform 1 0 23904 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_934
timestamp 1626908933
transform 1 0 23904 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_54
timestamp 1626908933
transform 1 0 24672 0 -1 27972
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_8
timestamp 1626908933
transform 1 0 24672 0 -1 27972
box -38 -49 2726 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_699
timestamp 1626908933
transform 1 0 26900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_51
timestamp 1626908933
transform 1 0 26900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_699
timestamp 1626908933
transform 1 0 26900 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_51
timestamp 1626908933
transform 1 0 26900 0 1 27306
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2300
timestamp 1626908933
transform 1 0 26928 0 1 27417
box -29 -23 29 23
use L1M1_PR  L1M1_PR_365
timestamp 1626908933
transform 1 0 26928 0 1 27417
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1944
timestamp 1626908933
transform 1 0 27360 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_953
timestamp 1626908933
transform 1 0 27360 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1109
timestamp 1626908933
transform 1 0 27552 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_118
timestamp 1626908933
transform 1 0 27552 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_838
timestamp 1626908933
transform 1 0 27648 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_116
timestamp 1626908933
transform 1 0 27648 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_414
timestamp 1626908933
transform 1 0 27456 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_57
timestamp 1626908933
transform 1 0 27456 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_36
timestamp 1626908933
transform -1 0 28896 0 -1 27972
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_11
timestamp 1626908933
transform -1 0 28896 0 -1 27972
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_675
timestamp 1626908933
transform 1 0 29300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_27
timestamp 1626908933
transform 1 0 29300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_675
timestamp 1626908933
transform 1 0 29300 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_27
timestamp 1626908933
transform 1 0 29300 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1108
timestamp 1626908933
transform 1 0 28896 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_117
timestamp 1626908933
transform 1 0 28896 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_804
timestamp 1626908933
transform 1 0 28992 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_82
timestamp 1626908933
transform 1 0 28992 0 -1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2308
timestamp 1626908933
transform 1 0 29904 0 1 27417
box -32 -32 32 32
use M1M2_PR  M1M2_PR_341
timestamp 1626908933
transform 1 0 29904 0 1 27417
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_663
timestamp 1626908933
transform 1 0 29760 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_62
timestamp 1626908933
transform 1 0 29760 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_624
timestamp 1626908933
transform 1 0 29952 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_26
timestamp 1626908933
transform 1 0 29952 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_758
timestamp 1626908933
transform 1 0 30336 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_36
timestamp 1626908933
transform 1 0 30336 0 -1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_602
timestamp 1626908933
transform 1 0 31104 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_4
timestamp 1626908933
transform 1 0 31104 0 -1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_116
timestamp 1626908933
transform 1 0 31488 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1107
timestamp 1626908933
transform 1 0 31488 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_56
timestamp 1626908933
transform 1 0 31680 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_413
timestamp 1626908933
transform 1 0 31680 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_954
timestamp 1626908933
transform 1 0 31584 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1945
timestamp 1626908933
transform 1 0 31584 0 -1 27972
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_3
timestamp 1626908933
transform 1 0 31700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_651
timestamp 1626908933
transform 1 0 31700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_3
timestamp 1626908933
transform 1 0 31700 0 1 27306
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_651
timestamp 1626908933
transform 1 0 31700 0 1 27306
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_579
timestamp 1626908933
transform 1 0 31776 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1180
timestamp 1626908933
transform 1 0 31776 0 -1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1946
timestamp 1626908933
transform 1 0 31968 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_955
timestamp 1626908933
transform 1 0 31968 0 -1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_55
timestamp 1626908933
transform 1 0 288 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_412
timestamp 1626908933
transform 1 0 288 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_580
timestamp 1626908933
transform 1 0 0 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1181
timestamp 1626908933
transform 1 0 0 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_956
timestamp 1626908933
transform 1 0 192 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1947
timestamp 1626908933
transform 1 0 192 0 1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1845
timestamp 1626908933
transform 1 0 48 0 1 27713
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3812
timestamp 1626908933
transform 1 0 48 0 1 27713
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_691
timestamp 1626908933
transform 1 0 768 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1413
timestamp 1626908933
transform 1 0 768 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_589
timestamp 1626908933
transform 1 0 384 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1187
timestamp 1626908933
transform 1 0 384 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_115
timestamp 1626908933
transform 1 0 1536 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1106
timestamp 1626908933
transform 1 0 1536 0 1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1122
timestamp 1626908933
transform 1 0 1488 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3089
timestamp 1626908933
transform 1 0 1488 0 1 27565
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_627
timestamp 1626908933
transform 1 0 1700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1275
timestamp 1626908933
transform 1 0 1700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_627
timestamp 1626908933
transform 1 0 1700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1275
timestamp 1626908933
transform 1 0 1700 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_558
timestamp 1626908933
transform 1 0 1632 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1156
timestamp 1626908933
transform 1 0 1632 0 1 27972
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3085
timestamp 1626908933
transform 1 0 2160 0 1 28083
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1118
timestamp 1626908933
transform 1 0 2160 0 1 28083
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1105
timestamp 1626908933
transform 1 0 2016 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_114
timestamp 1626908933
transform 1 0 2016 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1381
timestamp 1626908933
transform 1 0 2112 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_659
timestamp 1626908933
transform 1 0 2112 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_61
timestamp 1626908933
transform 1 0 2880 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_662
timestamp 1626908933
transform 1 0 2880 0 1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1194
timestamp 1626908933
transform 1 0 3024 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3129
timestamp 1626908933
transform 1 0 3024 0 1 27565
box -29 -23 29 23
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_41
timestamp 1626908933
transform 1 0 3072 0 1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_103
timestamp 1626908933
transform 1 0 3072 0 1 27972
box -38 -49 326 715
use L1M1_PR  L1M1_PR_1189
timestamp 1626908933
transform 1 0 3216 0 1 28083
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3124
timestamp 1626908933
transform 1 0 3216 0 1 28083
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_636
timestamp 1626908933
transform 1 0 3360 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1358
timestamp 1626908933
transform 1 0 3360 0 1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2170
timestamp 1626908933
transform 1 0 4272 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_203
timestamp 1626908933
transform 1 0 4272 0 1 27639
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1251
timestamp 1626908933
transform 1 0 4100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_603
timestamp 1626908933
transform 1 0 4100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1251
timestamp 1626908933
transform 1 0 4100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_603
timestamp 1626908933
transform 1 0 4100 0 1 27972
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3121
timestamp 1626908933
transform 1 0 4272 0 1 28231
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1186
timestamp 1626908933
transform 1 0 4272 0 1 28231
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1182
timestamp 1626908933
transform 1 0 4128 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_581
timestamp 1626908933
transform 1 0 4128 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_122
timestamp 1626908933
transform -1 0 4800 0 1 27972
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_53
timestamp 1626908933
transform -1 0 4800 0 1 27972
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1212
timestamp 1626908933
transform 1 0 4464 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3179
timestamp 1626908933
transform 1 0 4464 0 1 27565
box -32 -32 32 32
use L1M1_PR  L1M1_PR_223
timestamp 1626908933
transform 1 0 4560 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1284
timestamp 1626908933
transform 1 0 4464 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2158
timestamp 1626908933
transform 1 0 4560 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3219
timestamp 1626908933
transform 1 0 4464 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_316
timestamp 1626908933
transform 1 0 4656 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2251
timestamp 1626908933
transform 1 0 4656 0 1 27639
box -29 -23 29 23
use M1M2_PR  M1M2_PR_294
timestamp 1626908933
transform 1 0 4752 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2261
timestamp 1626908933
transform 1 0 4752 0 1 27639
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2250
timestamp 1626908933
transform 1 0 4848 0 1 28083
box -29 -23 29 23
use L1M1_PR  L1M1_PR_315
timestamp 1626908933
transform 1 0 4848 0 1 28083
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2260
timestamp 1626908933
transform 1 0 4752 0 1 28083
box -32 -32 32 32
use M1M2_PR  M1M2_PR_293
timestamp 1626908933
transform 1 0 4752 0 1 28083
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1183
timestamp 1626908933
transform 1 0 4800 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_582
timestamp 1626908933
transform 1 0 4800 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_54
timestamp 1626908933
transform 1 0 4992 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_411
timestamp 1626908933
transform 1 0 4992 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_113
timestamp 1626908933
transform 1 0 5088 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1104
timestamp 1626908933
transform 1 0 5088 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_597
timestamp 1626908933
transform 1 0 5184 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1319
timestamp 1626908933
transform 1 0 5184 0 1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_207
timestamp 1626908933
transform 1 0 5712 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1000
timestamp 1626908933
transform 1 0 6192 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2174
timestamp 1626908933
transform 1 0 5712 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2967
timestamp 1626908933
transform 1 0 6192 0 1 27861
box -32 -32 32 32
use L1M1_PR  L1M1_PR_227
timestamp 1626908933
transform 1 0 6192 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1064
timestamp 1626908933
transform 1 0 6288 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2162
timestamp 1626908933
transform 1 0 6192 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2999
timestamp 1626908933
transform 1 0 6288 0 1 27861
box -29 -23 29 23
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_25
timestamp 1626908933
transform 1 0 5952 0 1 27972
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_64
timestamp 1626908933
transform 1 0 5952 0 1 27972
box -38 -49 614 715
use M1M2_PR  M1M2_PR_996
timestamp 1626908933
transform 1 0 6672 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1163
timestamp 1626908933
transform 1 0 6384 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2963
timestamp 1626908933
transform 1 0 6672 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3130
timestamp 1626908933
transform 1 0 6384 0 1 27565
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1059
timestamp 1626908933
transform 1 0 6576 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2994
timestamp 1626908933
transform 1 0 6576 0 1 27861
box -29 -23 29 23
use M1M2_PR  M1M2_PR_995
timestamp 1626908933
transform 1 0 6672 0 1 28231
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2962
timestamp 1626908933
transform 1 0 6672 0 1 28231
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_579
timestamp 1626908933
transform 1 0 6500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1227
timestamp 1626908933
transform 1 0 6500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_579
timestamp 1626908933
transform 1 0 6500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1227
timestamp 1626908933
transform 1 0 6500 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_571
timestamp 1626908933
transform 1 0 6528 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1293
timestamp 1626908933
transform 1 0 6528 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_60
timestamp 1626908933
transform 1 0 7296 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_661
timestamp 1626908933
transform 1 0 7296 0 1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1684
timestamp 1626908933
transform 1 0 7632 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3619
timestamp 1626908933
transform 1 0 7632 0 1 27639
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1593
timestamp 1626908933
transform 1 0 7920 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3560
timestamp 1626908933
transform 1 0 7920 0 1 27639
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1716
timestamp 1626908933
transform 1 0 8016 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3651
timestamp 1626908933
transform 1 0 8016 0 1 27639
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_552
timestamp 1626908933
transform 1 0 7872 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1274
timestamp 1626908933
transform 1 0 7872 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_462
timestamp 1626908933
transform 1 0 7488 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1060
timestamp 1626908933
transform 1 0 7488 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_112
timestamp 1626908933
transform 1 0 8640 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1103
timestamp 1626908933
transform 1 0 8640 0 1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_199
timestamp 1626908933
transform 1 0 8688 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1629
timestamp 1626908933
transform 1 0 8304 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2166
timestamp 1626908933
transform 1 0 8688 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3596
timestamp 1626908933
transform 1 0 8304 0 1 27639
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_555
timestamp 1626908933
transform 1 0 8900 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1203
timestamp 1626908933
transform 1 0 8900 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_555
timestamp 1626908933
transform 1 0 8900 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1203
timestamp 1626908933
transform 1 0 8900 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_532
timestamp 1626908933
transform 1 0 8736 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1254
timestamp 1626908933
transform 1 0 8736 0 1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1093
timestamp 1626908933
transform 1 0 9264 0 1 28083
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3060
timestamp 1626908933
transform 1 0 9264 0 1 28083
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_44
timestamp 1626908933
transform 1 0 9504 0 1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_106
timestamp 1626908933
transform 1 0 9504 0 1 27972
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_583
timestamp 1626908933
transform 1 0 9792 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1184
timestamp 1626908933
transform 1 0 9792 0 1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1158
timestamp 1626908933
transform 1 0 9648 0 1 28083
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3093
timestamp 1626908933
transform 1 0 9648 0 1 28083
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_53
timestamp 1626908933
transform 1 0 9984 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_410
timestamp 1626908933
transform 1 0 9984 0 1 27972
box -38 -49 134 715
use L1M1_PR  L1M1_PR_219
timestamp 1626908933
transform 1 0 9936 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2154
timestamp 1626908933
transform 1 0 9936 0 1 27861
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1013
timestamp 1626908933
transform 1 0 10080 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_415
timestamp 1626908933
transform 1 0 10080 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1227
timestamp 1626908933
transform 1 0 10464 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_505
timestamp 1626908933
transform 1 0 10464 0 1 27972
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1179
timestamp 1626908933
transform 1 0 11300 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_531
timestamp 1626908933
transform 1 0 11300 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1179
timestamp 1626908933
transform 1 0 11300 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_531
timestamp 1626908933
transform 1 0 11300 0 1 27972
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3084
timestamp 1626908933
transform 1 0 11088 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1149
timestamp 1626908933
transform 1 0 11088 0 1 27861
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_660
timestamp 1626908933
transform 1 0 11232 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_59
timestamp 1626908933
transform 1 0 11232 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1102
timestamp 1626908933
transform 1 0 11424 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_111
timestamp 1626908933
transform 1 0 11424 0 1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1082
timestamp 1626908933
transform 1 0 12048 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3049
timestamp 1626908933
transform 1 0 12048 0 1 27861
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_477
timestamp 1626908933
transform 1 0 11520 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1199
timestamp 1626908933
transform 1 0 11520 0 1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1715
timestamp 1626908933
transform 1 0 13776 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3682
timestamp 1626908933
transform 1 0 13776 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_257
timestamp 1626908933
transform 1 0 12624 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2224
timestamp 1626908933
transform 1 0 12624 0 1 27861
box -32 -32 32 32
use L1M1_PR  L1M1_PR_280
timestamp 1626908933
transform 1 0 13488 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2215
timestamp 1626908933
transform 1 0 13488 0 1 27861
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_507
timestamp 1626908933
transform 1 0 13700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1155
timestamp 1626908933
transform 1 0 13700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_507
timestamp 1626908933
transform 1 0 13700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1155
timestamp 1626908933
transform 1 0 13700 0 1 27972
box -100 -49 100 49
use M1M2_PR  M1M2_PR_256
timestamp 1626908933
transform 1 0 12624 0 1 28083
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2223
timestamp 1626908933
transform 1 0 12624 0 1 28083
box -32 -32 32 32
use L1M1_PR  L1M1_PR_281
timestamp 1626908933
transform 1 0 12624 0 1 28083
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2216
timestamp 1626908933
transform 1 0 12624 0 1 28083
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_71
timestamp 1626908933
transform -1 0 14976 0 1 27972
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_25
timestamp 1626908933
transform -1 0 14976 0 1 27972
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1075
timestamp 1626908933
transform 1 0 13872 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3042
timestamp 1626908933
transform 1 0 13872 0 1 27639
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1141
timestamp 1626908933
transform 1 0 13872 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3076
timestamp 1626908933
transform 1 0 13872 0 1 27639
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1563
timestamp 1626908933
transform 1 0 14064 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3530
timestamp 1626908933
transform 1 0 14064 0 1 27861
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1652
timestamp 1626908933
transform 1 0 14064 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3587
timestamp 1626908933
transform 1 0 14064 0 1 27861
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1612
timestamp 1626908933
transform 1 0 14544 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3579
timestamp 1626908933
transform 1 0 14544 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1562
timestamp 1626908933
transform 1 0 14064 0 1 28231
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3529
timestamp 1626908933
transform 1 0 14064 0 1 28231
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3586
timestamp 1626908933
transform 1 0 14928 0 1 28231
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1651
timestamp 1626908933
transform 1 0 14928 0 1 28231
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1101
timestamp 1626908933
transform 1 0 15456 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_110
timestamp 1626908933
transform 1 0 15456 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_911
timestamp 1626908933
transform 1 0 15072 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_313
timestamp 1626908933
transform 1 0 15072 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_409
timestamp 1626908933
transform 1 0 14976 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_52
timestamp 1626908933
transform 1 0 14976 0 1 27972
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1131
timestamp 1626908933
transform 1 0 16100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_483
timestamp 1626908933
transform 1 0 16100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1131
timestamp 1626908933
transform 1 0 16100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_483
timestamp 1626908933
transform 1 0 16100 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1100
timestamp 1626908933
transform 1 0 16320 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_109
timestamp 1626908933
transform 1 0 16320 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1123
timestamp 1626908933
transform 1 0 15552 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_401
timestamp 1626908933
transform 1 0 15552 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_891
timestamp 1626908933
transform 1 0 16416 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_293
timestamp 1626908933
transform 1 0 16416 0 1 27972
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1606
timestamp 1626908933
transform 1 0 17040 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1607
timestamp 1626908933
transform 1 0 17040 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3573
timestamp 1626908933
transform 1 0 17040 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3574
timestamp 1626908933
transform 1 0 17040 0 1 27639
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1663
timestamp 1626908933
transform 1 0 17424 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1699
timestamp 1626908933
transform 1 0 17040 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3598
timestamp 1626908933
transform 1 0 17424 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3634
timestamp 1626908933
transform 1 0 17040 0 1 27639
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_374
timestamp 1626908933
transform 1 0 16800 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1096
timestamp 1626908933
transform 1 0 16800 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1099
timestamp 1626908933
transform 1 0 17568 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1098
timestamp 1626908933
transform 1 0 18048 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_108
timestamp 1626908933
transform 1 0 17568 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_107
timestamp 1626908933
transform 1 0 18048 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_856
timestamp 1626908933
transform 1 0 17664 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_258
timestamp 1626908933
transform 1 0 17664 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1069
timestamp 1626908933
transform 1 0 18144 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_347
timestamp 1626908933
transform 1 0 18144 0 1 27972
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_459
timestamp 1626908933
transform 1 0 18500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1107
timestamp 1626908933
transform 1 0 18500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_459
timestamp 1626908933
transform 1 0 18500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1107
timestamp 1626908933
transform 1 0 18500 0 1 27972
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1843
timestamp 1626908933
transform 1 0 18672 0 1 28231
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1844
timestamp 1626908933
transform 1 0 18672 0 1 27713
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3810
timestamp 1626908933
transform 1 0 18672 0 1 28231
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3811
timestamp 1626908933
transform 1 0 18672 0 1 27713
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_58
timestamp 1626908933
transform 1 0 18912 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_659
timestamp 1626908933
transform 1 0 18912 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_106
timestamp 1626908933
transform 1 0 19104 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1097
timestamp 1626908933
transform 1 0 19104 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1042
timestamp 1626908933
transform 1 0 19200 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_320
timestamp 1626908933
transform 1 0 19200 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1096
timestamp 1626908933
transform 1 0 20064 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_105
timestamp 1626908933
transform 1 0 20064 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_810
timestamp 1626908933
transform 1 0 20160 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_212
timestamp 1626908933
transform 1 0 20160 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_408
timestamp 1626908933
transform 1 0 19968 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_51
timestamp 1626908933
transform 1 0 19968 0 1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1430
timestamp 1626908933
transform 1 0 20976 0 1 27713
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3397
timestamp 1626908933
transform 1 0 20976 0 1 27713
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1822
timestamp 1626908933
transform 1 0 20592 0 1 28231
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3757
timestamp 1626908933
transform 1 0 20592 0 1 28231
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_435
timestamp 1626908933
transform 1 0 20900 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1083
timestamp 1626908933
transform 1 0 20900 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_435
timestamp 1626908933
transform 1 0 20900 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1083
timestamp 1626908933
transform 1 0 20900 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_0
timestamp 1626908933
transform 1 0 20544 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_6
timestamp 1626908933
transform 1 0 20544 0 1 27972
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3319
timestamp 1626908933
transform 1 0 21072 0 1 28083
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1384
timestamp 1626908933
transform 1 0 21072 0 1 28083
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3260
timestamp 1626908933
transform 1 0 21168 0 1 28083
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1293
timestamp 1626908933
transform 1 0 21168 0 1 28083
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1000
timestamp 1626908933
transform 1 0 21312 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_278
timestamp 1626908933
transform 1 0 21312 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_778
timestamp 1626908933
transform 1 0 22080 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_180
timestamp 1626908933
transform 1 0 22080 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1095
timestamp 1626908933
transform 1 0 22464 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_104
timestamp 1626908933
transform 1 0 22464 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_964
timestamp 1626908933
transform 1 0 22560 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_242
timestamp 1626908933
transform 1 0 22560 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_57
timestamp 1626908933
transform 1 0 23328 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_658
timestamp 1626908933
transform 1 0 23328 0 1 27972
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1498
timestamp 1626908933
transform 1 0 23280 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3433
timestamp 1626908933
transform 1 0 23280 0 1 27565
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_411
timestamp 1626908933
transform 1 0 23300 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1059
timestamp 1626908933
transform 1 0 23300 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_411
timestamp 1626908933
transform 1 0 23300 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1059
timestamp 1626908933
transform 1 0 23300 0 1 27972
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1512
timestamp 1626908933
transform 1 0 23472 0 1 27713
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3447
timestamp 1626908933
transform 1 0 23472 0 1 27713
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_153
timestamp 1626908933
transform 1 0 23520 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_751
timestamp 1626908933
transform 1 0 23520 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_933
timestamp 1626908933
transform 1 0 23904 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_211
timestamp 1626908933
transform 1 0 23904 0 1 27972
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3432
timestamp 1626908933
transform 1 0 24720 0 1 27565
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1497
timestamp 1626908933
transform 1 0 24720 0 1 27565
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1094
timestamp 1626908933
transform 1 0 24672 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_103
timestamp 1626908933
transform 1 0 24672 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1185
timestamp 1626908933
transform 1 0 24768 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_584
timestamp 1626908933
transform 1 0 24768 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_50
timestamp 1626908933
transform 1 0 24960 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_407
timestamp 1626908933
transform 1 0 24960 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_121
timestamp 1626908933
transform 1 0 25056 0 1 27972
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_719
timestamp 1626908933
transform 1 0 25056 0 1 27972
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1462
timestamp 1626908933
transform 1 0 25104 0 1 27639
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3397
timestamp 1626908933
transform 1 0 25104 0 1 27639
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1375
timestamp 1626908933
transform 1 0 25488 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3342
timestamp 1626908933
transform 1 0 25488 0 1 27639
box -32 -32 32 32
use L1M1_PR  L1M1_PR_369
timestamp 1626908933
transform 1 0 25776 0 1 28083
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2304
timestamp 1626908933
transform 1 0 25776 0 1 28083
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_387
timestamp 1626908933
transform 1 0 25700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1035
timestamp 1626908933
transform 1 0 25700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_387
timestamp 1626908933
transform 1 0 25700 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1035
timestamp 1626908933
transform 1 0 25700 0 1 27972
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1420
timestamp 1626908933
transform 1 0 26064 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3387
timestamp 1626908933
transform 1 0 26064 0 1 27639
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2346
timestamp 1626908933
transform 1 0 26544 0 1 27565
box -32 -32 32 32
use M1M2_PR  M1M2_PR_379
timestamp 1626908933
transform 1 0 26544 0 1 27565
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_49
timestamp 1626908933
transform -1 0 28128 0 1 27972
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_3
timestamp 1626908933
transform -1 0 28128 0 1 27972
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_346
timestamp 1626908933
transform 1 0 27696 0 1 28083
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2313
timestamp 1626908933
transform 1 0 27696 0 1 28083
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_363
timestamp 1626908933
transform 1 0 28100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1011
timestamp 1626908933
transform 1 0 28100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_363
timestamp 1626908933
transform 1 0 28100 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1011
timestamp 1626908933
transform 1 0 28100 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_56
timestamp 1626908933
transform 1 0 28128 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_657
timestamp 1626908933
transform 1 0 28128 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_102
timestamp 1626908933
transform 1 0 28320 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1093
timestamp 1626908933
transform 1 0 28320 0 1 27972
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1413
timestamp 1626908933
transform 1 0 28464 0 1 27861
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3380
timestamp 1626908933
transform 1 0 28464 0 1 27861
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_105
timestamp 1626908933
transform 1 0 28416 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_827
timestamp 1626908933
transform 1 0 28416 0 1 27972
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1354
timestamp 1626908933
transform 1 0 29136 0 1 27713
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3321
timestamp 1626908933
transform 1 0 29136 0 1 27713
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1438
timestamp 1626908933
transform 1 0 28848 0 1 27713
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1495
timestamp 1626908933
transform 1 0 28560 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1503
timestamp 1626908933
transform 1 0 28656 0 1 27713
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3373
timestamp 1626908933
transform 1 0 28848 0 1 27713
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3430
timestamp 1626908933
transform 1 0 28560 0 1 27861
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3438
timestamp 1626908933
transform 1 0 28656 0 1 27713
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_69
timestamp 1626908933
transform 1 0 29184 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_791
timestamp 1626908933
transform 1 0 29184 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_656
timestamp 1626908933
transform 1 0 30048 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_55
timestamp 1626908933
transform 1 0 30048 0 1 27972
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_406
timestamp 1626908933
transform 1 0 29952 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_49
timestamp 1626908933
transform 1 0 29952 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1092
timestamp 1626908933
transform 1 0 30240 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_101
timestamp 1626908933
transform 1 0 30240 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_757
timestamp 1626908933
transform 1 0 30336 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_35
timestamp 1626908933
transform 1 0 30336 0 1 27972
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_987
timestamp 1626908933
transform 1 0 30500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_339
timestamp 1626908933
transform 1 0 30500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_987
timestamp 1626908933
transform 1 0 30500 0 1 27972
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_339
timestamp 1626908933
transform 1 0 30500 0 1 27972
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1091
timestamp 1626908933
transform 1 0 31104 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_100
timestamp 1626908933
transform 1 0 31104 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_724
timestamp 1626908933
transform 1 0 31200 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_2
timestamp 1626908933
transform 1 0 31200 0 1 27972
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1948
timestamp 1626908933
transform 1 0 31968 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_957
timestamp 1626908933
transform 1 0 31968 0 1 27972
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_54
timestamp 1626908933
transform 1 0 0 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_655
timestamp 1626908933
transform 1 0 0 0 -1 29304
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1842
timestamp 1626908933
transform 1 0 144 0 1 28453
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3809
timestamp 1626908933
transform 1 0 144 0 1 28453
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_314
timestamp 1626908933
transform 1 0 500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_962
timestamp 1626908933
transform 1 0 500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_314
timestamp 1626908933
transform 1 0 500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_962
timestamp 1626908933
transform 1 0 500 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_702
timestamp 1626908933
transform 1 0 192 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1424
timestamp 1626908933
transform 1 0 192 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1090
timestamp 1626908933
transform 1 0 960 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_99
timestamp 1626908933
transform 1 0 960 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1162
timestamp 1626908933
transform 1 0 1056 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_564
timestamp 1626908933
transform 1 0 1056 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1390
timestamp 1626908933
transform 1 0 1440 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_668
timestamp 1626908933
transform 1 0 1440 0 -1 29304
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3084
timestamp 1626908933
transform 1 0 2160 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1117
timestamp 1626908933
transform 1 0 2160 0 1 28305
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1089
timestamp 1626908933
transform 1 0 2208 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_98
timestamp 1626908933
transform 1 0 2208 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1186
timestamp 1626908933
transform 1 0 2304 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_585
timestamp 1626908933
transform 1 0 2304 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_405
timestamp 1626908933
transform 1 0 2496 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_48
timestamp 1626908933
transform 1 0 2496 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1088
timestamp 1626908933
transform 1 0 2592 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_97
timestamp 1626908933
transform 1 0 2592 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1374
timestamp 1626908933
transform 1 0 2688 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_652
timestamp 1626908933
transform 1 0 2688 0 -1 29304
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3122
timestamp 1626908933
transform 1 0 3120 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1187
timestamp 1626908933
transform 1 0 3120 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3119
timestamp 1626908933
transform 1 0 3312 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1184
timestamp 1626908933
transform 1 0 3312 0 1 28305
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3080
timestamp 1626908933
transform 1 0 3312 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1113
timestamp 1626908933
transform 1 0 3312 0 1 28305
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_938
timestamp 1626908933
transform 1 0 2900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_290
timestamp 1626908933
transform 1 0 2900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_938
timestamp 1626908933
transform 1 0 2900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_290
timestamp 1626908933
transform 1 0 2900 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_532
timestamp 1626908933
transform 1 0 3456 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1130
timestamp 1626908933
transform 1 0 3456 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_654
timestamp 1626908933
transform 1 0 3840 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_53
timestamp 1626908933
transform 1 0 3840 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1346
timestamp 1626908933
transform 1 0 4032 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_624
timestamp 1626908933
transform 1 0 4032 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_96
timestamp 1626908933
transform 1 0 4800 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1087
timestamp 1626908933
transform 1 0 4800 0 -1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_266
timestamp 1626908933
transform 1 0 5300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_914
timestamp 1626908933
transform 1 0 5300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_266
timestamp 1626908933
transform 1 0 5300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_914
timestamp 1626908933
transform 1 0 5300 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_596
timestamp 1626908933
transform 1 0 5280 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1318
timestamp 1626908933
transform 1 0 5280 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_508
timestamp 1626908933
transform 1 0 4896 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1106
timestamp 1626908933
transform 1 0 4896 0 -1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2176
timestamp 1626908933
transform 1 0 5520 0 1 28379
box -32 -32 32 32
use M1M2_PR  M1M2_PR_209
timestamp 1626908933
transform 1 0 5520 0 1 28379
box -32 -32 32 32
use M1M2_PR  M1M2_PR_999
timestamp 1626908933
transform 1 0 6192 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1591
timestamp 1626908933
transform 1 0 6000 0 1 28527
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2966
timestamp 1626908933
transform 1 0 6192 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3558
timestamp 1626908933
transform 1 0 6000 0 1 28527
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1065
timestamp 1626908933
transform 1 0 6192 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1679
timestamp 1626908933
transform 1 0 6000 0 1 28527
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3000
timestamp 1626908933
transform 1 0 6192 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3614
timestamp 1626908933
transform 1 0 6000 0 1 28527
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_488
timestamp 1626908933
transform 1 0 6048 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1086
timestamp 1626908933
transform 1 0 6048 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_95
timestamp 1626908933
transform 1 0 6432 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1086
timestamp 1626908933
transform 1 0 6432 0 -1 29304
box -38 -49 134 715
use M1M2_PR  M1M2_PR_992
timestamp 1626908933
transform 1 0 6768 0 1 28971
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2959
timestamp 1626908933
transform 1 0 6768 0 1 28971
box -32 -32 32 32
use L1M1_PR  L1M1_PR_226
timestamp 1626908933
transform 1 0 6480 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1061
timestamp 1626908933
transform 1 0 6384 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2161
timestamp 1626908933
transform 1 0 6480 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2996
timestamp 1626908933
transform 1 0 6384 0 1 28305
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_570
timestamp 1626908933
transform 1 0 6528 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1292
timestamp 1626908933
transform 1 0 6528 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1949
timestamp 1626908933
transform 1 0 7392 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1085
timestamp 1626908933
transform 1 0 7296 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_958
timestamp 1626908933
transform 1 0 7392 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_94
timestamp 1626908933
transform 1 0 7296 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_404
timestamp 1626908933
transform 1 0 7488 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_47
timestamp 1626908933
transform 1 0 7488 0 -1 29304
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_890
timestamp 1626908933
transform 1 0 7700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_242
timestamp 1626908933
transform 1 0 7700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_890
timestamp 1626908933
transform 1 0 7700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_242
timestamp 1626908933
transform 1 0 7700 0 1 28638
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1592
timestamp 1626908933
transform 1 0 7920 0 1 28749
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3559
timestamp 1626908933
transform 1 0 7920 0 1 28749
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1683
timestamp 1626908933
transform 1 0 8016 0 1 28749
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3618
timestamp 1626908933
transform 1 0 8016 0 1 28749
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_461
timestamp 1626908933
transform 1 0 7584 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1059
timestamp 1626908933
transform 1 0 7584 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_24
timestamp 1626908933
transform 1 0 7968 0 -1 29304
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_63
timestamp 1626908933
transform 1 0 7968 0 -1 29304
box -38 -49 614 715
use L1M1_PR  L1M1_PR_2987
timestamp 1626908933
transform 1 0 8208 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1052
timestamp 1626908933
transform 1 0 8208 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2985
timestamp 1626908933
transform 1 0 8400 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2155
timestamp 1626908933
transform 1 0 8496 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1050
timestamp 1626908933
transform 1 0 8400 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_220
timestamp 1626908933
transform 1 0 8496 0 1 28971
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2955
timestamp 1626908933
transform 1 0 8304 0 1 28971
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2168
timestamp 1626908933
transform 1 0 8496 0 1 28971
box -32 -32 32 32
use M1M2_PR  M1M2_PR_988
timestamp 1626908933
transform 1 0 8304 0 1 28971
box -32 -32 32 32
use M1M2_PR  M1M2_PR_201
timestamp 1626908933
transform 1 0 8496 0 1 28971
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_653
timestamp 1626908933
transform 1 0 8544 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_52
timestamp 1626908933
transform 1 0 8544 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_531
timestamp 1626908933
transform 1 0 9120 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1253
timestamp 1626908933
transform 1 0 9120 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_443
timestamp 1626908933
transform 1 0 8736 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1041
timestamp 1626908933
transform 1 0 8736 0 -1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1087
timestamp 1626908933
transform 1 0 9456 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3054
timestamp 1626908933
transform 1 0 9456 0 1 28305
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1154
timestamp 1626908933
transform 1 0 9552 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3089
timestamp 1626908933
transform 1 0 9552 0 1 28305
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_51
timestamp 1626908933
transform 1 0 9888 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_652
timestamp 1626908933
transform 1 0 9888 0 -1 29304
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1083
timestamp 1626908933
transform 1 0 9840 0 1 28971
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1084
timestamp 1626908933
transform 1 0 9840 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3050
timestamp 1626908933
transform 1 0 9840 0 1 28971
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3051
timestamp 1626908933
transform 1 0 9840 0 1 28305
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1152
timestamp 1626908933
transform 1 0 9744 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3087
timestamp 1626908933
transform 1 0 9744 0 1 28305
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_866
timestamp 1626908933
transform 1 0 10100 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_218
timestamp 1626908933
transform 1 0 10100 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_866
timestamp 1626908933
transform 1 0 10100 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_218
timestamp 1626908933
transform 1 0 10100 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1012
timestamp 1626908933
transform 1 0 10080 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_414
timestamp 1626908933
transform 1 0 10080 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1226
timestamp 1626908933
transform 1 0 10464 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_504
timestamp 1626908933
transform 1 0 10464 0 -1 29304
box -38 -49 806 715
use M1M2_PR  M1M2_PR_262
timestamp 1626908933
transform 1 0 11472 0 1 29045
box -32 -32 32 32
use M1M2_PR  M1M2_PR_265
timestamp 1626908933
transform 1 0 11856 0 1 28749
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2229
timestamp 1626908933
transform 1 0 11472 0 1 29045
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2232
timestamp 1626908933
transform 1 0 11856 0 1 28749
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1150
timestamp 1626908933
transform 1 0 11856 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3085
timestamp 1626908933
transform 1 0 11856 0 1 28971
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_391
timestamp 1626908933
transform 1 0 11232 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_989
timestamp 1626908933
transform 1 0 11232 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_33
timestamp 1626908933
transform 1 0 11616 0 -1 29304
box -38 -49 614 715
use sky130_fd_sc_hs__o21a_1  sky130_fd_sc_hs__o21a_1_72
timestamp 1626908933
transform 1 0 11616 0 -1 29304
box -38 -49 614 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_586
timestamp 1626908933
transform 1 0 12192 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1187
timestamp 1626908933
transform 1 0 12192 0 -1 29304
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1081
timestamp 1626908933
transform 1 0 12048 0 1 28897
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3048
timestamp 1626908933
transform 1 0 12048 0 1 28897
box -32 -32 32 32
use L1M1_PR  L1M1_PR_287
timestamp 1626908933
transform 1 0 12240 0 1 28749
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1148
timestamp 1626908933
transform 1 0 12048 0 1 28897
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2222
timestamp 1626908933
transform 1 0 12240 0 1 28749
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3083
timestamp 1626908933
transform 1 0 12048 0 1 28897
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_46
timestamp 1626908933
transform 1 0 12480 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_403
timestamp 1626908933
transform 1 0 12480 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_959
timestamp 1626908933
transform 1 0 12384 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1950
timestamp 1626908933
transform 1 0 12384 0 -1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_194
timestamp 1626908933
transform 1 0 12500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_842
timestamp 1626908933
transform 1 0 12500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_194
timestamp 1626908933
transform 1 0 12500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_842
timestamp 1626908933
transform 1 0 12500 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_357
timestamp 1626908933
transform 1 0 12576 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_955
timestamp 1626908933
transform 1 0 12576 0 -1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3686
timestamp 1626908933
transform 1 0 13488 0 1 28379
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1719
timestamp 1626908933
transform 1 0 13488 0 1 28379
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1175
timestamp 1626908933
transform 1 0 12960 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_453
timestamp 1626908933
transform 1 0 12960 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_49
timestamp 1626908933
transform -1 0 14208 0 -1 29304
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_118
timestamp 1626908933
transform -1 0 14208 0 -1 29304
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_93
timestamp 1626908933
transform 1 0 14208 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1084
timestamp 1626908933
transform 1 0 14208 0 -1 29304
box -38 -49 134 715
use M1M2_PR  M1M2_PR_261
timestamp 1626908933
transform 1 0 13968 0 1 29045
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1074
timestamp 1626908933
transform 1 0 13968 0 1 28749
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2228
timestamp 1626908933
transform 1 0 13968 0 1 29045
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3041
timestamp 1626908933
transform 1 0 13968 0 1 28749
box -32 -32 32 32
use L1M1_PR  L1M1_PR_284
timestamp 1626908933
transform 1 0 13872 0 1 28971
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2219
timestamp 1626908933
transform 1 0 13872 0 1 28971
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1611
timestamp 1626908933
transform 1 0 14544 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3578
timestamp 1626908933
transform 1 0 14544 0 1 28305
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1704
timestamp 1626908933
transform 1 0 14544 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3639
timestamp 1626908933
transform 1 0 14544 0 1 28305
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_426
timestamp 1626908933
transform 1 0 14304 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1148
timestamp 1626908933
transform 1 0 14304 0 -1 29304
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_818
timestamp 1626908933
transform 1 0 14900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_170
timestamp 1626908933
transform 1 0 14900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_818
timestamp 1626908933
transform 1 0 14900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_170
timestamp 1626908933
transform 1 0 14900 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1083
timestamp 1626908933
transform 1 0 15456 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_92
timestamp 1626908933
transform 1 0 15456 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_910
timestamp 1626908933
transform 1 0 15072 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_312
timestamp 1626908933
transform 1 0 15072 0 -1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3040
timestamp 1626908933
transform 1 0 16272 0 1 28749
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1073
timestamp 1626908933
transform 1 0 16272 0 1 28749
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1951
timestamp 1626908933
transform 1 0 16320 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_960
timestamp 1626908933
transform 1 0 16320 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1122
timestamp 1626908933
transform 1 0 15552 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_400
timestamp 1626908933
transform 1 0 15552 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_107
timestamp 1626908933
transform -1 0 16704 0 -1 29304
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_45
timestamp 1626908933
transform -1 0 16704 0 -1 29304
box -38 -49 326 715
use L1M1_PR  L1M1_PR_3082
timestamp 1626908933
transform 1 0 16464 0 1 28897
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3074
timestamp 1626908933
transform 1 0 16368 0 1 28749
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1147
timestamp 1626908933
transform 1 0 16464 0 1 28897
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1139
timestamp 1626908933
transform 1 0 16368 0 1 28749
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_794
timestamp 1626908933
transform 1 0 17300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_146
timestamp 1626908933
transform 1 0 17300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_794
timestamp 1626908933
transform 1 0 17300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_146
timestamp 1626908933
transform 1 0 17300 0 1 28638
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3047
timestamp 1626908933
transform 1 0 16656 0 1 28897
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1080
timestamp 1626908933
transform 1 0 16656 0 1 28897
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_44
timestamp 1626908933
transform 1 0 16704 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_21
timestamp 1626908933
transform 1 0 16704 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_45
timestamp 1626908933
transform 1 0 17472 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_402
timestamp 1626908933
transform 1 0 17472 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_91
timestamp 1626908933
transform 1 0 17568 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1082
timestamp 1626908933
transform 1 0 17568 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_90
timestamp 1626908933
transform 1 0 18048 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1081
timestamp 1626908933
transform 1 0 18048 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_346
timestamp 1626908933
transform 1 0 18144 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1068
timestamp 1626908933
transform 1 0 18144 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_257
timestamp 1626908933
transform 1 0 17664 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_855
timestamp 1626908933
transform 1 0 17664 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1080
timestamp 1626908933
transform 1 0 18912 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_89
timestamp 1626908933
transform 1 0 18912 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_833
timestamp 1626908933
transform 1 0 19008 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_235
timestamp 1626908933
transform 1 0 19008 0 -1 29304
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_770
timestamp 1626908933
transform 1 0 19700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_122
timestamp 1626908933
transform 1 0 19700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_770
timestamp 1626908933
transform 1 0 19700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_122
timestamp 1626908933
transform 1 0 19700 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1079
timestamp 1626908933
transform 1 0 20160 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_88
timestamp 1626908933
transform 1 0 20160 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1041
timestamp 1626908933
transform 1 0 19392 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_319
timestamp 1626908933
transform 1 0 19392 0 -1 29304
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3322
timestamp 1626908933
transform 1 0 20880 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1387
timestamp 1626908933
transform 1 0 20880 0 1 28305
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3271
timestamp 1626908933
transform 1 0 20688 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1304
timestamp 1626908933
transform 1 0 20688 0 1 28305
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_809
timestamp 1626908933
transform 1 0 20256 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_211
timestamp 1626908933
transform 1 0 20256 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1016
timestamp 1626908933
transform 1 0 20640 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_294
timestamp 1626908933
transform 1 0 20640 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1078
timestamp 1626908933
transform 1 0 21600 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_87
timestamp 1626908933
transform 1 0 21600 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_651
timestamp 1626908933
transform 1 0 21408 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_50
timestamp 1626908933
transform 1 0 21408 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_987
timestamp 1626908933
transform 1 0 21696 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_265
timestamp 1626908933
transform 1 0 21696 0 -1 29304
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_746
timestamp 1626908933
transform 1 0 22100 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_98
timestamp 1626908933
transform 1 0 22100 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_746
timestamp 1626908933
transform 1 0 22100 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_98
timestamp 1626908933
transform 1 0 22100 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_963
timestamp 1626908933
transform 1 0 22560 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_241
timestamp 1626908933
transform 1 0 22560 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_401
timestamp 1626908933
transform 1 0 22464 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_44
timestamp 1626908933
transform 1 0 22464 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_650
timestamp 1626908933
transform 1 0 23328 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_49
timestamp 1626908933
transform 1 0 23328 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_750
timestamp 1626908933
transform 1 0 23520 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_152
timestamp 1626908933
transform 1 0 23520 0 -1 29304
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_722
timestamp 1626908933
transform 1 0 24500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_74
timestamp 1626908933
transform 1 0 24500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_722
timestamp 1626908933
transform 1 0 24500 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_74
timestamp 1626908933
transform 1 0 24500 0 1 28638
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3808
timestamp 1626908933
transform 1 0 24048 0 1 28453
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1841
timestamp 1626908933
transform 1 0 24048 0 1 28453
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_932
timestamp 1626908933
transform 1 0 23904 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_210
timestamp 1626908933
transform 1 0 23904 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1077
timestamp 1626908933
transform 1 0 24672 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_86
timestamp 1626908933
transform 1 0 24672 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_726
timestamp 1626908933
transform 1 0 24768 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_128
timestamp 1626908933
transform 1 0 24768 0 -1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3341
timestamp 1626908933
transform 1 0 25488 0 1 28305
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1374
timestamp 1626908933
transform 1 0 25488 0 1 28305
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_898
timestamp 1626908933
transform 1 0 25152 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_176
timestamp 1626908933
transform 1 0 25152 0 -1 29304
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2345
timestamp 1626908933
transform 1 0 26544 0 1 28379
box -32 -32 32 32
use M1M2_PR  M1M2_PR_378
timestamp 1626908933
transform 1 0 26544 0 1 28379
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_649
timestamp 1626908933
transform 1 0 25920 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_48
timestamp 1626908933
transform 1 0 25920 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_698
timestamp 1626908933
transform 1 0 26112 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_100
timestamp 1626908933
transform 1 0 26112 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_870
timestamp 1626908933
transform 1 0 26496 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_148
timestamp 1626908933
transform 1 0 26496 0 -1 29304
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_698
timestamp 1626908933
transform 1 0 26900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_50
timestamp 1626908933
transform 1 0 26900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_698
timestamp 1626908933
transform 1 0 26900 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_50
timestamp 1626908933
transform 1 0 26900 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1952
timestamp 1626908933
transform 1 0 27360 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1076
timestamp 1626908933
transform 1 0 27264 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_961
timestamp 1626908933
transform 1 0 27360 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_85
timestamp 1626908933
transform 1 0 27264 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_648
timestamp 1626908933
transform 1 0 27552 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_47
timestamp 1626908933
transform 1 0 27552 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_400
timestamp 1626908933
transform 1 0 27456 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_43
timestamp 1626908933
transform 1 0 27456 0 -1 29304
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3431
timestamp 1626908933
transform 1 0 28080 0 1 28379
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3390
timestamp 1626908933
transform 1 0 27696 0 1 28305
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1496
timestamp 1626908933
transform 1 0 28080 0 1 28379
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1455
timestamp 1626908933
transform 1 0 27696 0 1 28305
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3379
timestamp 1626908933
transform 1 0 28464 0 1 28379
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1412
timestamp 1626908933
transform 1 0 28464 0 1 28379
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_837
timestamp 1626908933
transform 1 0 27744 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_115
timestamp 1626908933
transform 1 0 27744 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_84
timestamp 1626908933
transform 1 0 28896 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1075
timestamp 1626908933
transform 1 0 28896 0 -1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_26
timestamp 1626908933
transform 1 0 29300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_674
timestamp 1626908933
transform 1 0 29300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_26
timestamp 1626908933
transform 1 0 29300 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_674
timestamp 1626908933
transform 1 0 29300 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_81
timestamp 1626908933
transform 1 0 28992 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_803
timestamp 1626908933
transform 1 0 28992 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_55
timestamp 1626908933
transform 1 0 28512 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_653
timestamp 1626908933
transform 1 0 28512 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_647
timestamp 1626908933
transform 1 0 29760 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_46
timestamp 1626908933
transform 1 0 29760 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_623
timestamp 1626908933
transform 1 0 29952 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_25
timestamp 1626908933
transform 1 0 29952 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_756
timestamp 1626908933
transform 1 0 30336 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_34
timestamp 1626908933
transform 1 0 30336 0 -1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_601
timestamp 1626908933
transform 1 0 31104 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_3
timestamp 1626908933
transform 1 0 31104 0 -1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_83
timestamp 1626908933
transform 1 0 31488 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1074
timestamp 1626908933
transform 1 0 31488 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_42
timestamp 1626908933
transform 1 0 31680 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_399
timestamp 1626908933
transform 1 0 31680 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_962
timestamp 1626908933
transform 1 0 31584 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1953
timestamp 1626908933
transform 1 0 31584 0 -1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_2
timestamp 1626908933
transform 1 0 31700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_650
timestamp 1626908933
transform 1 0 31700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_2
timestamp 1626908933
transform 1 0 31700 0 1 28638
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_650
timestamp 1626908933
transform 1 0 31700 0 1 28638
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_587
timestamp 1626908933
transform 1 0 31776 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1188
timestamp 1626908933
transform 1 0 31776 0 -1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1954
timestamp 1626908933
transform 1 0 31968 0 -1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_963
timestamp 1626908933
transform 1 0 31968 0 -1 29304
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3806
timestamp 1626908933
transform 1 0 48 0 1 29489
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1839
timestamp 1626908933
transform 1 0 48 0 1 29489
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1955
timestamp 1626908933
transform 1 0 192 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_964
timestamp 1626908933
transform 1 0 192 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1189
timestamp 1626908933
transform 1 0 0 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_588
timestamp 1626908933
transform 1 0 0 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_398
timestamp 1626908933
transform 1 0 288 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_41
timestamp 1626908933
transform 1 0 288 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1186
timestamp 1626908933
transform 1 0 384 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_588
timestamp 1626908933
transform 1 0 384 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_690
timestamp 1626908933
transform 1 0 768 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1412
timestamp 1626908933
transform 1 0 768 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_557
timestamp 1626908933
transform 1 0 1536 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1155
timestamp 1626908933
transform 1 0 1536 0 1 29304
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_626
timestamp 1626908933
transform 1 0 1700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1274
timestamp 1626908933
transform 1 0 1700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_626
timestamp 1626908933
transform 1 0 1700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1274
timestamp 1626908933
transform 1 0 1700 0 1 29304
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1119
timestamp 1626908933
transform 1 0 1968 0 1 29563
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3086
timestamp 1626908933
transform 1 0 1968 0 1 29563
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1191
timestamp 1626908933
transform 1 0 1968 0 1 29563
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3126
timestamp 1626908933
transform 1 0 1968 0 1 29563
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1116
timestamp 1626908933
transform 1 0 2160 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3083
timestamp 1626908933
transform 1 0 2160 0 1 29637
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1188
timestamp 1626908933
transform 1 0 2160 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3123
timestamp 1626908933
transform 1 0 2160 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1185
timestamp 1626908933
transform 1 0 2256 0 1 29563
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3120
timestamp 1626908933
transform 1 0 2256 0 1 29563
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_112
timestamp 1626908933
transform -1 0 2304 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_50
timestamp 1626908933
transform -1 0 2304 0 1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1641
timestamp 1626908933
transform 1 0 2736 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3608
timestamp 1626908933
transform 1 0 2736 0 1 29637
box -32 -32 32 32
use L1M1_PR  L1M1_PR_229
timestamp 1626908933
transform 1 0 2736 0 1 29785
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2164
timestamp 1626908933
transform 1 0 2736 0 1 29785
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_80
timestamp 1626908933
transform -1 0 4992 0 1 29304
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_34
timestamp 1626908933
transform -1 0 4992 0 1 29304
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_3605
timestamp 1626908933
transform 1 0 3408 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3134
timestamp 1626908933
transform 1 0 3120 0 1 29711
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3079
timestamp 1626908933
transform 1 0 3312 0 1 29563
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1638
timestamp 1626908933
transform 1 0 3408 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1167
timestamp 1626908933
transform 1 0 3120 0 1 29711
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1112
timestamp 1626908933
transform 1 0 3312 0 1 29563
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1250
timestamp 1626908933
transform 1 0 4100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_602
timestamp 1626908933
transform 1 0 4100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1250
timestamp 1626908933
transform 1 0 4100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_602
timestamp 1626908933
transform 1 0 4100 0 1 29304
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1722
timestamp 1626908933
transform 1 0 4560 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3657
timestamp 1626908933
transform 1 0 4560 0 1 29637
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_40
timestamp 1626908933
transform 1 0 4992 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_397
timestamp 1626908933
transform 1 0 4992 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_45
timestamp 1626908933
transform 1 0 5088 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_646
timestamp 1626908933
transform 1 0 5088 0 1 29304
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1680
timestamp 1626908933
transform 1 0 4944 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3615
timestamp 1626908933
transform 1 0 4944 0 1 29637
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_595
timestamp 1626908933
transform 1 0 5280 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1317
timestamp 1626908933
transform 1 0 5280 0 1 29304
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2175
timestamp 1626908933
transform 1 0 5520 0 1 29785
box -32 -32 32 32
use M1M2_PR  M1M2_PR_208
timestamp 1626908933
transform 1 0 5520 0 1 29785
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_487
timestamp 1626908933
transform 1 0 6048 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1085
timestamp 1626908933
transform 1 0 6048 0 1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1590
timestamp 1626908933
transform 1 0 6000 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3557
timestamp 1626908933
transform 1 0 6000 0 1 29637
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_82
timestamp 1626908933
transform 1 0 6432 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1073
timestamp 1626908933
transform 1 0 6432 0 1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_578
timestamp 1626908933
transform 1 0 6500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1226
timestamp 1626908933
transform 1 0 6500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_578
timestamp 1626908933
transform 1 0 6500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1226
timestamp 1626908933
transform 1 0 6500 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_569
timestamp 1626908933
transform 1 0 6528 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1291
timestamp 1626908933
transform 1 0 6528 0 1 29304
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1631
timestamp 1626908933
transform 1 0 7536 0 1 29563
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3598
timestamp 1626908933
transform 1 0 7536 0 1 29563
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1718
timestamp 1626908933
transform 1 0 7728 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3653
timestamp 1626908933
transform 1 0 7728 0 1 29637
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1595
timestamp 1626908933
transform 1 0 7440 0 1 29711
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3562
timestamp 1626908933
transform 1 0 7440 0 1 29711
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1686
timestamp 1626908933
transform 1 0 7344 0 1 29711
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3621
timestamp 1626908933
transform 1 0 7344 0 1 29711
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1740
timestamp 1626908933
transform 1 0 8112 0 1 29711
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3707
timestamp 1626908933
transform 1 0 8112 0 1 29711
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_89
timestamp 1626908933
transform 1 0 7296 0 1 29304
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_43
timestamp 1626908933
transform 1 0 7296 0 1 29304
box -38 -49 2726 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1202
timestamp 1626908933
transform 1 0 8900 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_554
timestamp 1626908933
transform 1 0 8900 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1202
timestamp 1626908933
transform 1 0 8900 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_554
timestamp 1626908933
transform 1 0 8900 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_396
timestamp 1626908933
transform 1 0 9984 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_39
timestamp 1626908933
transform 1 0 9984 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1011
timestamp 1626908933
transform 1 0 10080 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_413
timestamp 1626908933
transform 1 0 10080 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1225
timestamp 1626908933
transform 1 0 10464 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_503
timestamp 1626908933
transform 1 0 10464 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_390
timestamp 1626908933
transform 1 0 11328 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_988
timestamp 1626908933
transform 1 0 11328 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_81
timestamp 1626908933
transform 1 0 11232 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1072
timestamp 1626908933
transform 1 0 11232 0 1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_530
timestamp 1626908933
transform 1 0 11300 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1178
timestamp 1626908933
transform 1 0 11300 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_530
timestamp 1626908933
transform 1 0 11300 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1178
timestamp 1626908933
transform 1 0 11300 0 1 29304
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3583
timestamp 1626908933
transform 1 0 11664 0 1 29193
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1648
timestamp 1626908933
transform 1 0 11664 0 1 29193
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2231
timestamp 1626908933
transform 1 0 11856 0 1 29785
box -32 -32 32 32
use M1M2_PR  M1M2_PR_264
timestamp 1626908933
transform 1 0 11856 0 1 29785
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1956
timestamp 1626908933
transform 1 0 11808 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1071
timestamp 1626908933
transform 1 0 11712 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_965
timestamp 1626908933
transform 1 0 11808 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_80
timestamp 1626908933
transform 1 0 11712 0 1 29304
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3582
timestamp 1626908933
transform 1 0 11952 0 1 29563
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1647
timestamp 1626908933
transform 1 0 11952 0 1 29563
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3526
timestamp 1626908933
transform 1 0 11952 0 1 29193
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3525
timestamp 1626908933
transform 1 0 11952 0 1 29563
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1559
timestamp 1626908933
transform 1 0 11952 0 1 29193
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1558
timestamp 1626908933
transform 1 0 11952 0 1 29563
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1621
timestamp 1626908933
transform 1 0 12336 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3588
timestamp 1626908933
transform 1 0 12336 0 1 29637
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1708
timestamp 1626908933
transform 1 0 12336 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3643
timestamp 1626908933
transform 1 0 12336 0 1 29637
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1154
timestamp 1626908933
transform 1 0 13700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_506
timestamp 1626908933
transform 1 0 13700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1154
timestamp 1626908933
transform 1 0 13700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_506
timestamp 1626908933
transform 1 0 13700 0 1 29304
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3685
timestamp 1626908933
transform 1 0 13488 0 1 29711
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1718
timestamp 1626908933
transform 1 0 13488 0 1 29711
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_74
timestamp 1626908933
transform 1 0 11904 0 1 29304
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_28
timestamp 1626908933
transform 1 0 11904 0 1 29304
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_3080
timestamp 1626908933
transform 1 0 14064 0 1 29119
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2221
timestamp 1626908933
transform 1 0 14160 0 1 29785
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1145
timestamp 1626908933
transform 1 0 14064 0 1 29119
box -29 -23 29 23
use L1M1_PR  L1M1_PR_286
timestamp 1626908933
transform 1 0 14160 0 1 29785
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3577
timestamp 1626908933
transform 1 0 14544 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1610
timestamp 1626908933
transform 1 0 14544 0 1 29637
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_925
timestamp 1626908933
transform 1 0 14592 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_327
timestamp 1626908933
transform 1 0 14592 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1070
timestamp 1626908933
transform 1 0 15456 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_79
timestamp 1626908933
transform 1 0 15456 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_909
timestamp 1626908933
transform 1 0 15072 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_311
timestamp 1626908933
transform 1 0 15072 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_395
timestamp 1626908933
transform 1 0 14976 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_38
timestamp 1626908933
transform 1 0 14976 0 1 29304
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1072
timestamp 1626908933
transform 1 0 16272 0 1 29415
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3039
timestamp 1626908933
transform 1 0 16272 0 1 29415
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1140
timestamp 1626908933
transform 1 0 16272 0 1 29415
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3075
timestamp 1626908933
transform 1 0 16272 0 1 29415
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_482
timestamp 1626908933
transform 1 0 16100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1130
timestamp 1626908933
transform 1 0 16100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_482
timestamp 1626908933
transform 1 0 16100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1130
timestamp 1626908933
transform 1 0 16100 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_399
timestamp 1626908933
transform 1 0 15552 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1121
timestamp 1626908933
transform 1 0 15552 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_46
timestamp 1626908933
transform 1 0 16320 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_108
timestamp 1626908933
transform 1 0 16320 0 1 29304
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3079
timestamp 1626908933
transform 1 0 16464 0 1 29637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1144
timestamp 1626908933
transform 1 0 16464 0 1 29637
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3045
timestamp 1626908933
transform 1 0 16464 0 1 29119
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3044
timestamp 1626908933
transform 1 0 16464 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1078
timestamp 1626908933
transform 1 0 16464 0 1 29119
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1077
timestamp 1626908933
transform 1 0 16464 0 1 29637
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_78
timestamp 1626908933
transform 1 0 16704 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1069
timestamp 1626908933
transform 1 0 16704 0 1 29304
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1079
timestamp 1626908933
transform 1 0 16656 0 1 29563
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3046
timestamp 1626908933
transform 1 0 16656 0 1 29563
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1143
timestamp 1626908933
transform 1 0 16752 0 1 29119
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1146
timestamp 1626908933
transform 1 0 16656 0 1 29563
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3078
timestamp 1626908933
transform 1 0 16752 0 1 29119
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3081
timestamp 1626908933
transform 1 0 16656 0 1 29563
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_373
timestamp 1626908933
transform 1 0 16800 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1095
timestamp 1626908933
transform 1 0 16800 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1068
timestamp 1626908933
transform 1 0 17568 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1067
timestamp 1626908933
transform 1 0 18048 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_77
timestamp 1626908933
transform 1 0 17568 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_76
timestamp 1626908933
transform 1 0 18048 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_854
timestamp 1626908933
transform 1 0 17664 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_256
timestamp 1626908933
transform 1 0 17664 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1067
timestamp 1626908933
transform 1 0 18144 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_345
timestamp 1626908933
transform 1 0 18144 0 1 29304
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1106
timestamp 1626908933
transform 1 0 18500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_458
timestamp 1626908933
transform 1 0 18500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1106
timestamp 1626908933
transform 1 0 18500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_458
timestamp 1626908933
transform 1 0 18500 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1066
timestamp 1626908933
transform 1 0 19104 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_75
timestamp 1626908933
transform 1 0 19104 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_645
timestamp 1626908933
transform 1 0 18912 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_44
timestamp 1626908933
transform 1 0 18912 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1040
timestamp 1626908933
transform 1 0 19200 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_318
timestamp 1626908933
transform 1 0 19200 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1026
timestamp 1626908933
transform 1 0 20064 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_304
timestamp 1626908933
transform 1 0 20064 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_394
timestamp 1626908933
transform 1 0 19968 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_37
timestamp 1626908933
transform 1 0 19968 0 1 29304
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1082
timestamp 1626908933
transform 1 0 20900 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_434
timestamp 1626908933
transform 1 0 20900 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1082
timestamp 1626908933
transform 1 0 20900 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_434
timestamp 1626908933
transform 1 0 20900 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1065
timestamp 1626908933
transform 1 0 20832 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_74
timestamp 1626908933
transform 1 0 20832 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_798
timestamp 1626908933
transform 1 0 20928 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_200
timestamp 1626908933
transform 1 0 20928 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_999
timestamp 1626908933
transform 1 0 21312 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_277
timestamp 1626908933
transform 1 0 21312 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_777
timestamp 1626908933
transform 1 0 22080 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_179
timestamp 1626908933
transform 1 0 22080 0 1 29304
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3804
timestamp 1626908933
transform 1 0 22320 0 1 29489
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1837
timestamp 1626908933
transform 1 0 22320 0 1 29489
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1064
timestamp 1626908933
transform 1 0 22464 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_73
timestamp 1626908933
transform 1 0 22464 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_962
timestamp 1626908933
transform 1 0 22560 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_240
timestamp 1626908933
transform 1 0 22560 0 1 29304
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1058
timestamp 1626908933
transform 1 0 23300 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_410
timestamp 1626908933
transform 1 0 23300 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1058
timestamp 1626908933
transform 1 0 23300 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_410
timestamp 1626908933
transform 1 0 23300 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_644
timestamp 1626908933
transform 1 0 23328 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_43
timestamp 1626908933
transform 1 0 23328 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_749
timestamp 1626908933
transform 1 0 23520 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_151
timestamp 1626908933
transform 1 0 23520 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_931
timestamp 1626908933
transform 1 0 23904 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_209
timestamp 1626908933
transform 1 0 23904 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1957
timestamp 1626908933
transform 1 0 24864 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_966
timestamp 1626908933
transform 1 0 24864 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1190
timestamp 1626908933
transform 1 0 24672 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_589
timestamp 1626908933
transform 1 0 24672 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_36
timestamp 1626908933
transform 1 0 24960 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_393
timestamp 1626908933
transform 1 0 24960 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_72
timestamp 1626908933
transform 1 0 25056 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1063
timestamp 1626908933
transform 1 0 25056 0 1 29304
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_386
timestamp 1626908933
transform 1 0 25700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1034
timestamp 1626908933
transform 1 0 25700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_386
timestamp 1626908933
transform 1 0 25700 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1034
timestamp 1626908933
transform 1 0 25700 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_175
timestamp 1626908933
transform 1 0 25152 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_897
timestamp 1626908933
transform 1 0 25152 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_643
timestamp 1626908933
transform 1 0 25920 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_42
timestamp 1626908933
transform 1 0 25920 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_697
timestamp 1626908933
transform 1 0 26112 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_99
timestamp 1626908933
transform 1 0 26112 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_869
timestamp 1626908933
transform 1 0 26496 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_147
timestamp 1626908933
transform 1 0 26496 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1062
timestamp 1626908933
transform 1 0 27264 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_71
timestamp 1626908933
transform 1 0 27264 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_678
timestamp 1626908933
transform 1 0 27360 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_80
timestamp 1626908933
transform 1 0 27360 0 1 29304
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1010
timestamp 1626908933
transform 1 0 28100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_362
timestamp 1626908933
transform 1 0 28100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1010
timestamp 1626908933
transform 1 0 28100 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_362
timestamp 1626908933
transform 1 0 28100 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_836
timestamp 1626908933
transform 1 0 27744 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_114
timestamp 1626908933
transform 1 0 27744 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1061
timestamp 1626908933
transform 1 0 28896 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_70
timestamp 1626908933
transform 1 0 28896 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_652
timestamp 1626908933
transform 1 0 28512 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_54
timestamp 1626908933
transform 1 0 28512 0 1 29304
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_802
timestamp 1626908933
transform 1 0 28992 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_80
timestamp 1626908933
transform 1 0 28992 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1958
timestamp 1626908933
transform 1 0 29856 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1060
timestamp 1626908933
transform 1 0 29760 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_967
timestamp 1626908933
transform 1 0 29856 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_69
timestamp 1626908933
transform 1 0 29760 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_642
timestamp 1626908933
transform 1 0 30048 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_41
timestamp 1626908933
transform 1 0 30048 0 1 29304
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_392
timestamp 1626908933
transform 1 0 29952 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_35
timestamp 1626908933
transform 1 0 29952 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1059
timestamp 1626908933
transform 1 0 30240 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_68
timestamp 1626908933
transform 1 0 30240 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_755
timestamp 1626908933
transform 1 0 30336 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_33
timestamp 1626908933
transform 1 0 30336 0 1 29304
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_338
timestamp 1626908933
transform 1 0 30500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_986
timestamp 1626908933
transform 1 0 30500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_338
timestamp 1626908933
transform 1 0 30500 0 1 29304
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_986
timestamp 1626908933
transform 1 0 30500 0 1 29304
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_67
timestamp 1626908933
transform 1 0 31104 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1058
timestamp 1626908933
transform 1 0 31104 0 1 29304
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1826
timestamp 1626908933
transform 1 0 30960 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3793
timestamp 1626908933
transform 1 0 30960 0 1 29637
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1
timestamp 1626908933
transform 1 0 31200 0 1 29304
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_723
timestamp 1626908933
transform 1 0 31200 0 1 29304
box -38 -49 806 715
use M1M2_PR  M1M2_PR_3791
timestamp 1626908933
transform 1 0 31920 0 1 29637
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1824
timestamp 1626908933
transform 1 0 31920 0 1 29637
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1959
timestamp 1626908933
transform 1 0 31968 0 1 29304
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_968
timestamp 1626908933
transform 1 0 31968 0 1 29304
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_961
timestamp 1626908933
transform 1 0 500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_313
timestamp 1626908933
transform 1 0 500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_961
timestamp 1626908933
transform 1 0 500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_313
timestamp 1626908933
transform 1 0 500 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_641
timestamp 1626908933
transform 1 0 0 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_40
timestamp 1626908933
transform 1 0 0 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1423
timestamp 1626908933
transform 1 0 192 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_701
timestamp 1626908933
transform 1 0 192 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1057
timestamp 1626908933
transform 1 0 960 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_66
timestamp 1626908933
transform 1 0 960 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1161
timestamp 1626908933
transform 1 0 1056 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_563
timestamp 1626908933
transform 1 0 1056 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1389
timestamp 1626908933
transform 1 0 1440 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_667
timestamp 1626908933
transform 1 0 1440 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_65
timestamp 1626908933
transform 1 0 2208 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1056
timestamp 1626908933
transform 1 0 2208 0 -1 30636
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1544
timestamp 1626908933
transform 1 0 2064 0 1 30229
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1545
timestamp 1626908933
transform 1 0 2064 0 1 29859
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3511
timestamp 1626908933
transform 1 0 2064 0 1 30229
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3512
timestamp 1626908933
transform 1 0 2064 0 1 29859
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1634
timestamp 1626908933
transform 1 0 1968 0 1 29859
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3569
timestamp 1626908933
transform 1 0 1968 0 1 29859
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_34
timestamp 1626908933
transform 1 0 2496 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_391
timestamp 1626908933
transform 1 0 2496 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_590
timestamp 1626908933
transform 1 0 2304 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1191
timestamp 1626908933
transform 1 0 2304 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1192
timestamp 1626908933
transform 1 0 2592 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_591
timestamp 1626908933
transform 1 0 2592 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_969
timestamp 1626908933
transform 1 0 2784 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1960
timestamp 1626908933
transform 1 0 2784 0 -1 30636
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1633
timestamp 1626908933
transform 1 0 2928 0 1 30229
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3568
timestamp 1626908933
transform 1 0 2928 0 1 30229
box -29 -23 29 23
use fine_freq_track_VIA0  fine_freq_track_VIA0_289
timestamp 1626908933
transform 1 0 2900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_937
timestamp 1626908933
transform 1 0 2900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_289
timestamp 1626908933
transform 1 0 2900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_937
timestamp 1626908933
transform 1 0 2900 0 1 29970
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1166
timestamp 1626908933
transform 1 0 3120 0 1 30229
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3133
timestamp 1626908933
transform 1 0 3120 0 1 30229
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1640
timestamp 1626908933
transform 1 0 3312 0 1 30303
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3607
timestamp 1626908933
transform 1 0 3312 0 1 30303
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1724
timestamp 1626908933
transform 1 0 3312 0 1 30303
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3659
timestamp 1626908933
transform 1 0 3312 0 1 30303
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_913
timestamp 1626908933
transform 1 0 5300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_265
timestamp 1626908933
transform 1 0 5300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_913
timestamp 1626908933
transform 1 0 5300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_265
timestamp 1626908933
transform 1 0 5300 0 1 29970
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2249
timestamp 1626908933
transform 1 0 5136 0 1 30081
box -29 -23 29 23
use L1M1_PR  L1M1_PR_314
timestamp 1626908933
transform 1 0 5136 0 1 30081
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2259
timestamp 1626908933
transform 1 0 4752 0 1 30081
box -32 -32 32 32
use M1M2_PR  M1M2_PR_292
timestamp 1626908933
transform 1 0 4752 0 1 30081
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_81
timestamp 1626908933
transform 1 0 2880 0 -1 30636
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_35
timestamp 1626908933
transform 1 0 2880 0 -1 30636
box -38 -49 2726 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1096
timestamp 1626908933
transform 1 0 5568 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_498
timestamp 1626908933
transform 1 0 5568 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1309
timestamp 1626908933
transform 1 0 5952 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_587
timestamp 1626908933
transform 1 0 5952 0 -1 30636
box -38 -49 806 715
use M1M2_PR  M1M2_PR_2958
timestamp 1626908933
transform 1 0 6768 0 1 30451
box -32 -32 32 32
use M1M2_PR  M1M2_PR_991
timestamp 1626908933
transform 1 0 6768 0 1 30451
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1287
timestamp 1626908933
transform 1 0 6720 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_565
timestamp 1626908933
transform 1 0 6720 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_33
timestamp 1626908933
transform 1 0 7488 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_390
timestamp 1626908933
transform 1 0 7488 0 -1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_241
timestamp 1626908933
transform 1 0 7700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_889
timestamp 1626908933
transform 1 0 7700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_241
timestamp 1626908933
transform 1 0 7700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_889
timestamp 1626908933
transform 1 0 7700 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_592
timestamp 1626908933
transform 1 0 7968 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1193
timestamp 1626908933
transform 1 0 7968 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_460
timestamp 1626908933
transform 1 0 7584 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1058
timestamp 1626908933
transform 1 0 7584 0 -1 30636
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2986
timestamp 1626908933
transform 1 0 8208 0 1 30451
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2157
timestamp 1626908933
transform 1 0 8112 0 1 30081
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1051
timestamp 1626908933
transform 1 0 8208 0 1 30451
box -29 -23 29 23
use L1M1_PR  L1M1_PR_222
timestamp 1626908933
transform 1 0 8112 0 1 30081
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_111
timestamp 1626908933
transform -1 0 8448 0 -1 30636
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_50
timestamp 1626908933
transform -1 0 8448 0 -1 30636
box -38 -49 326 715
use M1M2_PR  M1M2_PR_200
timestamp 1626908933
transform 1 0 8496 0 1 30081
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2167
timestamp 1626908933
transform 1 0 8496 0 1 30081
box -32 -32 32 32
use M1M2_PR  M1M2_PR_984
timestamp 1626908933
transform 1 0 8688 0 1 30525
box -32 -32 32 32
use M1M2_PR  M1M2_PR_987
timestamp 1626908933
transform 1 0 8304 0 1 30377
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2951
timestamp 1626908933
transform 1 0 8688 0 1 30525
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2954
timestamp 1626908933
transform 1 0 8304 0 1 30377
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1049
timestamp 1626908933
transform 1 0 8400 0 1 30377
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2984
timestamp 1626908933
transform 1 0 8400 0 1 30377
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_545
timestamp 1626908933
transform 1 0 8448 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1267
timestamp 1626908933
transform 1 0 8448 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_593
timestamp 1626908933
transform 1 0 9216 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1194
timestamp 1626908933
transform 1 0 9216 0 -1 30636
box -38 -49 230 715
use L1M1_PR  L1M1_PR_218
timestamp 1626908933
transform 1 0 9552 0 1 29859
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1044
timestamp 1626908933
transform 1 0 9552 0 1 30525
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2153
timestamp 1626908933
transform 1 0 9552 0 1 29859
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2979
timestamp 1626908933
transform 1 0 9552 0 1 30525
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_39
timestamp 1626908933
transform 1 0 9888 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_640
timestamp 1626908933
transform 1 0 9888 0 -1 30636
box -38 -49 230 715
use M1M2_PR  M1M2_PR_196
timestamp 1626908933
transform 1 0 9744 0 1 30303
box -32 -32 32 32
use M1M2_PR  M1M2_PR_197
timestamp 1626908933
transform 1 0 9744 0 1 29859
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2163
timestamp 1626908933
transform 1 0 9744 0 1 30303
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2164
timestamp 1626908933
transform 1 0 9744 0 1 29859
box -32 -32 32 32
use L1M1_PR  L1M1_PR_216
timestamp 1626908933
transform 1 0 9744 0 1 30303
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2151
timestamp 1626908933
transform 1 0 9744 0 1 30303
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_109
timestamp 1626908933
transform 1 0 9408 0 -1 30636
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_40
timestamp 1626908933
transform 1 0 9408 0 -1 30636
box -38 -49 518 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_865
timestamp 1626908933
transform 1 0 10100 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_217
timestamp 1626908933
transform 1 0 10100 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_865
timestamp 1626908933
transform 1 0 10100 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_217
timestamp 1626908933
transform 1 0 10100 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1010
timestamp 1626908933
transform 1 0 10080 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_412
timestamp 1626908933
transform 1 0 10080 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1224
timestamp 1626908933
transform 1 0 10464 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_502
timestamp 1626908933
transform 1 0 10464 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1055
timestamp 1626908933
transform 1 0 11232 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_64
timestamp 1626908933
transform 1 0 11232 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_987
timestamp 1626908933
transform 1 0 11328 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_389
timestamp 1626908933
transform 1 0 11328 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1198
timestamp 1626908933
transform 1 0 11712 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_476
timestamp 1626908933
transform 1 0 11712 0 -1 30636
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_841
timestamp 1626908933
transform 1 0 12500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_193
timestamp 1626908933
transform 1 0 12500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_841
timestamp 1626908933
transform 1 0 12500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_193
timestamp 1626908933
transform 1 0 12500 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_954
timestamp 1626908933
transform 1 0 12576 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_356
timestamp 1626908933
transform 1 0 12576 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_389
timestamp 1626908933
transform 1 0 12480 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_32
timestamp 1626908933
transform 1 0 12480 0 -1 30636
box -38 -49 134 715
use M1M2_PR  M1M2_PR_3684
timestamp 1626908933
transform 1 0 13488 0 1 30229
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1717
timestamp 1626908933
transform 1 0 13488 0 1 30229
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1174
timestamp 1626908933
transform 1 0 12960 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_452
timestamp 1626908933
transform 1 0 12960 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_639
timestamp 1626908933
transform 1 0 13728 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_38
timestamp 1626908933
transform 1 0 13728 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_63
timestamp 1626908933
transform 1 0 13920 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1054
timestamp 1626908933
transform 1 0 13920 0 -1 30636
box -38 -49 134 715
use M1M2_PR  M1M2_PR_260
timestamp 1626908933
transform 1 0 13968 0 1 30081
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2227
timestamp 1626908933
transform 1 0 13968 0 1 30081
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_169
timestamp 1626908933
transform 1 0 14900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_817
timestamp 1626908933
transform 1 0 14900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_169
timestamp 1626908933
transform 1 0 14900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_817
timestamp 1626908933
transform 1 0 14900 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_425
timestamp 1626908933
transform 1 0 14016 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1147
timestamp 1626908933
transform 1 0 14016 0 -1 30636
box -38 -49 806 715
use L1M1_PR  L1M1_PR_2218
timestamp 1626908933
transform 1 0 15216 0 1 30081
box -29 -23 29 23
use L1M1_PR  L1M1_PR_283
timestamp 1626908933
transform 1 0 15216 0 1 30081
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_84
timestamp 1626908933
transform -1 0 17472 0 -1 30636
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_38
timestamp 1626908933
transform -1 0 17472 0 -1 30636
box -38 -49 2726 715
use L1M1_PR  L1M1_PR_1650
timestamp 1626908933
transform 1 0 16656 0 1 29859
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3585
timestamp 1626908933
transform 1 0 16656 0 1 29859
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1561
timestamp 1626908933
transform 1 0 17136 0 1 29859
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3528
timestamp 1626908933
transform 1 0 17136 0 1 29859
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_145
timestamp 1626908933
transform 1 0 17300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_793
timestamp 1626908933
transform 1 0 17300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_145
timestamp 1626908933
transform 1 0 17300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_793
timestamp 1626908933
transform 1 0 17300 0 1 29970
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1560
timestamp 1626908933
transform 1 0 17136 0 1 30303
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1605
timestamp 1626908933
transform 1 0 17040 0 1 30303
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3527
timestamp 1626908933
transform 1 0 17136 0 1 30303
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3572
timestamp 1626908933
transform 1 0 17040 0 1 30303
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1698
timestamp 1626908933
transform 1 0 17040 0 1 30303
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3633
timestamp 1626908933
transform 1 0 17040 0 1 30303
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1649
timestamp 1626908933
transform 1 0 17424 0 1 30303
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3584
timestamp 1626908933
transform 1 0 17424 0 1 30303
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_31
timestamp 1626908933
transform 1 0 17472 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_388
timestamp 1626908933
transform 1 0 17472 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_62
timestamp 1626908933
transform 1 0 17568 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1053
timestamp 1626908933
transform 1 0 17568 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_61
timestamp 1626908933
transform 1 0 18048 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1052
timestamp 1626908933
transform 1 0 18048 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_344
timestamp 1626908933
transform 1 0 18144 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1066
timestamp 1626908933
transform 1 0 18144 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_255
timestamp 1626908933
transform 1 0 17664 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_853
timestamp 1626908933
transform 1 0 17664 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1051
timestamp 1626908933
transform 1 0 18912 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_60
timestamp 1626908933
transform 1 0 18912 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_832
timestamp 1626908933
transform 1 0 19008 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_234
timestamp 1626908933
transform 1 0 19008 0 -1 30636
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_769
timestamp 1626908933
transform 1 0 19700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_121
timestamp 1626908933
transform 1 0 19700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_769
timestamp 1626908933
transform 1 0 19700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_121
timestamp 1626908933
transform 1 0 19700 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1050
timestamp 1626908933
transform 1 0 20160 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_59
timestamp 1626908933
transform 1 0 20160 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1039
timestamp 1626908933
transform 1 0 19392 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_317
timestamp 1626908933
transform 1 0 19392 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_808
timestamp 1626908933
transform 1 0 20256 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_210
timestamp 1626908933
transform 1 0 20256 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1015
timestamp 1626908933
transform 1 0 20640 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_293
timestamp 1626908933
transform 1 0 20640 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1049
timestamp 1626908933
transform 1 0 21600 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_58
timestamp 1626908933
transform 1 0 21600 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_638
timestamp 1626908933
transform 1 0 21408 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_37
timestamp 1626908933
transform 1 0 21408 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_986
timestamp 1626908933
transform 1 0 21696 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_264
timestamp 1626908933
transform 1 0 21696 0 -1 30636
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_745
timestamp 1626908933
transform 1 0 22100 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_97
timestamp 1626908933
transform 1 0 22100 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_745
timestamp 1626908933
transform 1 0 22100 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_97
timestamp 1626908933
transform 1 0 22100 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_961
timestamp 1626908933
transform 1 0 22560 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_239
timestamp 1626908933
transform 1 0 22560 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_387
timestamp 1626908933
transform 1 0 22464 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_30
timestamp 1626908933
transform 1 0 22464 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_637
timestamp 1626908933
transform 1 0 23328 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_36
timestamp 1626908933
transform 1 0 23328 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_748
timestamp 1626908933
transform 1 0 23520 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_150
timestamp 1626908933
transform 1 0 23520 0 -1 30636
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_721
timestamp 1626908933
transform 1 0 24500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_73
timestamp 1626908933
transform 1 0 24500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_721
timestamp 1626908933
transform 1 0 24500 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_73
timestamp 1626908933
transform 1 0 24500 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_930
timestamp 1626908933
transform 1 0 23904 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_208
timestamp 1626908933
transform 1 0 23904 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1048
timestamp 1626908933
transform 1 0 24672 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_57
timestamp 1626908933
transform 1 0 24672 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_725
timestamp 1626908933
transform 1 0 24768 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_127
timestamp 1626908933
transform 1 0 24768 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_896
timestamp 1626908933
transform 1 0 25152 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_174
timestamp 1626908933
transform 1 0 25152 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_636
timestamp 1626908933
transform 1 0 25920 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_35
timestamp 1626908933
transform 1 0 25920 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_696
timestamp 1626908933
transform 1 0 26112 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_98
timestamp 1626908933
transform 1 0 26112 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_868
timestamp 1626908933
transform 1 0 26496 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_146
timestamp 1626908933
transform 1 0 26496 0 -1 30636
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_697
timestamp 1626908933
transform 1 0 26900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_49
timestamp 1626908933
transform 1 0 26900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_697
timestamp 1626908933
transform 1 0 26900 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_49
timestamp 1626908933
transform 1 0 26900 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1961
timestamp 1626908933
transform 1 0 27360 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1047
timestamp 1626908933
transform 1 0 27264 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_970
timestamp 1626908933
transform 1 0 27360 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_56
timestamp 1626908933
transform 1 0 27264 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_635
timestamp 1626908933
transform 1 0 27552 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_34
timestamp 1626908933
transform 1 0 27552 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_386
timestamp 1626908933
transform 1 0 27456 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_29
timestamp 1626908933
transform 1 0 27456 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_835
timestamp 1626908933
transform 1 0 27744 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_113
timestamp 1626908933
transform 1 0 27744 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_55
timestamp 1626908933
transform 1 0 28896 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1046
timestamp 1626908933
transform 1 0 28896 0 -1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_25
timestamp 1626908933
transform 1 0 29300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_673
timestamp 1626908933
transform 1 0 29300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_25
timestamp 1626908933
transform 1 0 29300 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_673
timestamp 1626908933
transform 1 0 29300 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_79
timestamp 1626908933
transform 1 0 28992 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_801
timestamp 1626908933
transform 1 0 28992 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_53
timestamp 1626908933
transform 1 0 28512 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_651
timestamp 1626908933
transform 1 0 28512 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_634
timestamp 1626908933
transform 1 0 29760 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_33
timestamp 1626908933
transform 1 0 29760 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_622
timestamp 1626908933
transform 1 0 29952 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_24
timestamp 1626908933
transform 1 0 29952 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_754
timestamp 1626908933
transform 1 0 30336 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_32
timestamp 1626908933
transform 1 0 30336 0 -1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_600
timestamp 1626908933
transform 1 0 31104 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_2
timestamp 1626908933
transform 1 0 31104 0 -1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_54
timestamp 1626908933
transform 1 0 31488 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1045
timestamp 1626908933
transform 1 0 31488 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_28
timestamp 1626908933
transform 1 0 31680 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_385
timestamp 1626908933
transform 1 0 31680 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_971
timestamp 1626908933
transform 1 0 31584 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1962
timestamp 1626908933
transform 1 0 31584 0 -1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_1
timestamp 1626908933
transform 1 0 31700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_649
timestamp 1626908933
transform 1 0 31700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1
timestamp 1626908933
transform 1 0 31700 0 1 29970
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_649
timestamp 1626908933
transform 1 0 31700 0 1 29970
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_594
timestamp 1626908933
transform 1 0 31776 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1195
timestamp 1626908933
transform 1 0 31776 0 -1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1963
timestamp 1626908933
transform 1 0 31968 0 -1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_972
timestamp 1626908933
transform 1 0 31968 0 -1 30636
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1836
timestamp 1626908933
transform 1 0 48 0 1 31117
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3803
timestamp 1626908933
transform 1 0 48 0 1 31117
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_27
timestamp 1626908933
transform 1 0 288 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_384
timestamp 1626908933
transform 1 0 288 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_973
timestamp 1626908933
transform 1 0 192 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1964
timestamp 1626908933
transform 1 0 192 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_26
timestamp 1626908933
transform 1 0 0 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_595
timestamp 1626908933
transform 1 0 0 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_627
timestamp 1626908933
transform 1 0 0 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1196
timestamp 1626908933
transform 1 0 0 0 1 30636
box -38 -49 230 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_960
timestamp 1626908933
transform 1 0 500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_312
timestamp 1626908933
transform 1 0 500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_960
timestamp 1626908933
transform 1 0 500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_312
timestamp 1626908933
transform 1 0 500 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1185
timestamp 1626908933
transform 1 0 384 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_587
timestamp 1626908933
transform 1 0 384 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_562
timestamp 1626908933
transform 1 0 1056 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1160
timestamp 1626908933
transform 1 0 1056 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_35
timestamp 1626908933
transform 1 0 960 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1026
timestamp 1626908933
transform 1 0 960 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_689
timestamp 1626908933
transform 1 0 768 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_700
timestamp 1626908933
transform 1 0 192 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1411
timestamp 1626908933
transform 1 0 768 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1422
timestamp 1626908933
transform 1 0 192 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1965
timestamp 1626908933
transform 1 0 1536 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_974
timestamp 1626908933
transform 1 0 1536 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1273
timestamp 1626908933
transform 1 0 1700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_625
timestamp 1626908933
transform 1 0 1700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1273
timestamp 1626908933
transform 1 0 1700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_625
timestamp 1626908933
transform 1 0 1700 0 1 30636
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2160
timestamp 1626908933
transform 1 0 2064 0 1 31191
box -29 -23 29 23
use L1M1_PR  L1M1_PR_225
timestamp 1626908933
transform 1 0 2064 0 1 31191
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2173
timestamp 1626908933
transform 1 0 2064 0 1 31191
box -32 -32 32 32
use M1M2_PR  M1M2_PR_206
timestamp 1626908933
transform 1 0 2064 0 1 31191
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_20
timestamp 1626908933
transform 1 0 2496 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_377
timestamp 1626908933
transform 1 0 2496 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_597
timestamp 1626908933
transform 1 0 2304 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1198
timestamp 1626908933
transform 1 0 2304 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_33
timestamp 1626908933
transform 1 0 2592 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_34
timestamp 1626908933
transform 1 0 2208 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1024
timestamp 1626908933
transform 1 0 2592 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1025
timestamp 1626908933
transform 1 0 2208 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_651
timestamp 1626908933
transform 1 0 2688 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_666
timestamp 1626908933
transform 1 0 1440 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1373
timestamp 1626908933
transform 1 0 2688 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1388
timestamp 1626908933
transform 1 0 1440 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_72
timestamp 1626908933
transform -1 0 4320 0 1 30636
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_26
timestamp 1626908933
transform -1 0 4320 0 1 30636
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_1165
timestamp 1626908933
transform 1 0 3120 0 1 31043
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1639
timestamp 1626908933
transform 1 0 3312 0 1 30969
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3132
timestamp 1626908933
transform 1 0 3120 0 1 31043
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3606
timestamp 1626908933
transform 1 0 3312 0 1 30969
box -32 -32 32 32
use fine_freq_track_VIA0  fine_freq_track_VIA0_288
timestamp 1626908933
transform 1 0 2900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_936
timestamp 1626908933
transform 1 0 2900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_288
timestamp 1626908933
transform 1 0 2900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_936
timestamp 1626908933
transform 1 0 2900 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_531
timestamp 1626908933
transform 1 0 3456 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1129
timestamp 1626908933
transform 1 0 3456 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_32
timestamp 1626908933
transform 1 0 3840 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1023
timestamp 1626908933
transform 1 0 3840 0 -1 31968
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1723
timestamp 1626908933
transform 1 0 3888 0 1 30969
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3658
timestamp 1626908933
transform 1 0 3888 0 1 30969
box -29 -23 29 23
use fine_freq_track_VIA1  fine_freq_track_VIA1_1249
timestamp 1626908933
transform 1 0 4100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_601
timestamp 1626908933
transform 1 0 4100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1249
timestamp 1626908933
transform 1 0 4100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_601
timestamp 1626908933
transform 1 0 4100 0 1 30636
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3617
timestamp 1626908933
transform 1 0 4272 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1682
timestamp 1626908933
transform 1 0 4272 0 1 30895
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_633
timestamp 1626908933
transform 1 0 4320 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_626
timestamp 1626908933
transform 1 0 4416 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_32
timestamp 1626908933
transform 1 0 4320 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_25
timestamp 1626908933
transform 1 0 4416 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_110
timestamp 1626908933
transform -1 0 4416 0 -1 31968
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_41
timestamp 1626908933
transform -1 0 4416 0 -1 31968
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_53
timestamp 1626908933
transform 1 0 4512 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1044
timestamp 1626908933
transform 1 0 4512 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_26
timestamp 1626908933
transform 1 0 4992 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_383
timestamp 1626908933
transform 1 0 4992 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_31
timestamp 1626908933
transform 1 0 5088 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_632
timestamp 1626908933
transform 1 0 5088 0 1 30636
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_264
timestamp 1626908933
transform 1 0 5300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_912
timestamp 1626908933
transform 1 0 5300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_264
timestamp 1626908933
transform 1 0 5300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_912
timestamp 1626908933
transform 1 0 5300 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_594
timestamp 1626908933
transform 1 0 5280 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_614
timestamp 1626908933
transform 1 0 4608 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1316
timestamp 1626908933
transform 1 0 5280 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1336
timestamp 1626908933
transform 1 0 4608 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_514
timestamp 1626908933
transform 1 0 4608 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1112
timestamp 1626908933
transform 1 0 4608 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_625
timestamp 1626908933
transform 1 0 5376 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_24
timestamp 1626908933
transform 1 0 5376 0 -1 31968
box -38 -49 230 715
use M1M2_PR  M1M2_PR_2965
timestamp 1626908933
transform 1 0 6288 0 1 30895
box -32 -32 32 32
use M1M2_PR  M1M2_PR_998
timestamp 1626908933
transform 1 0 6288 0 1 30895
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1022
timestamp 1626908933
transform 1 0 5568 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_31
timestamp 1626908933
transform 1 0 5568 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1084
timestamp 1626908933
transform 1 0 6048 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_486
timestamp 1626908933
transform 1 0 6048 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1308
timestamp 1626908933
transform 1 0 5664 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_586
timestamp 1626908933
transform 1 0 5664 0 -1 31968
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_577
timestamp 1626908933
transform 1 0 6500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1225
timestamp 1626908933
transform 1 0 6500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_577
timestamp 1626908933
transform 1 0 6500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1225
timestamp 1626908933
transform 1 0 6500 0 1 30636
box -100 -49 100 49
use L1M1_PR  L1M1_PR_1681
timestamp 1626908933
transform 1 0 6576 0 1 30821
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3616
timestamp 1626908933
transform 1 0 6576 0 1 30821
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1060
timestamp 1626908933
transform 1 0 6480 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2995
timestamp 1626908933
transform 1 0 6480 0 1 30895
box -29 -23 29 23
use M1M2_PR  M1M2_PR_990
timestamp 1626908933
transform 1 0 6768 0 1 30895
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2957
timestamp 1626908933
transform 1 0 6768 0 1 30895
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1054
timestamp 1626908933
transform 1 0 6768 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2989
timestamp 1626908933
transform 1 0 6768 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2990
timestamp 1626908933
transform 1 0 6672 0 1 30969
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1055
timestamp 1626908933
transform 1 0 6672 0 1 30969
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2961
timestamp 1626908933
transform 1 0 6576 0 1 30969
box -32 -32 32 32
use M1M2_PR  M1M2_PR_994
timestamp 1626908933
transform 1 0 6576 0 1 30969
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_115
timestamp 1626908933
transform 1 0 6432 0 -1 31968
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_53
timestamp 1626908933
transform 1 0 6432 0 -1 31968
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_564
timestamp 1626908933
transform 1 0 7200 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1286
timestamp 1626908933
transform 1 0 7200 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_477
timestamp 1626908933
transform 1 0 6816 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1075
timestamp 1626908933
transform 1 0 6816 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_22
timestamp 1626908933
transform 1 0 6720 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_45
timestamp 1626908933
transform 1 0 6720 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_38
timestamp 1626908933
transform -1 0 6816 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_100
timestamp 1626908933
transform -1 0 6816 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_888
timestamp 1626908933
transform 1 0 7700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_240
timestamp 1626908933
transform 1 0 7700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_888
timestamp 1626908933
transform 1 0 7700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_240
timestamp 1626908933
transform 1 0 7700 0 1 31302
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3561
timestamp 1626908933
transform 1 0 7440 0 1 30747
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1594
timestamp 1626908933
transform 1 0 7440 0 1 30747
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_376
timestamp 1626908933
transform 1 0 7488 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_19
timestamp 1626908933
transform 1 0 7488 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_624
timestamp 1626908933
transform 1 0 7584 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_23
timestamp 1626908933
transform 1 0 7584 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_551
timestamp 1626908933
transform 1 0 7776 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1273
timestamp 1626908933
transform 1 0 7776 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_457
timestamp 1626908933
transform 1 0 7968 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1055
timestamp 1626908933
transform 1 0 7968 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_52
timestamp 1626908933
transform 1 0 8352 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1043
timestamp 1626908933
transform 1 0 8352 0 1 30636
box -38 -49 134 715
use M1M2_PR  M1M2_PR_983
timestamp 1626908933
transform 1 0 8688 0 1 30969
box -32 -32 32 32
use M1M2_PR  M1M2_PR_985
timestamp 1626908933
transform 1 0 8400 0 1 30895
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2950
timestamp 1626908933
transform 1 0 8688 0 1 30969
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2952
timestamp 1626908933
transform 1 0 8400 0 1 30895
box -32 -32 32 32
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_54
timestamp 1626908933
transform 1 0 8544 0 -1 31968
box -38 -49 326 715
use sky130_fd_sc_hs__nor2_1  sky130_fd_sc_hs__nor2_1_116
timestamp 1626908933
transform 1 0 8544 0 -1 31968
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_22
timestamp 1626908933
transform 1 0 8832 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_623
timestamp 1626908933
transform 1 0 8832 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_30
timestamp 1626908933
transform 1 0 9024 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1021
timestamp 1626908933
transform 1 0 9024 0 -1 31968
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_553
timestamp 1626908933
transform 1 0 8900 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1201
timestamp 1626908933
transform 1 0 8900 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_553
timestamp 1626908933
transform 1 0 8900 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1201
timestamp 1626908933
transform 1 0 8900 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_530
timestamp 1626908933
transform 1 0 9120 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_544
timestamp 1626908933
transform 1 0 8448 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1252
timestamp 1626908933
transform 1 0 9120 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1266
timestamp 1626908933
transform 1 0 8448 0 1 30636
box -38 -49 806 715
use L1M1_PR  L1M1_PR_3620
timestamp 1626908933
transform 1 0 9360 0 1 30747
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1685
timestamp 1626908933
transform 1 0 9360 0 1 30747
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2982
timestamp 1626908933
transform 1 0 9264 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1047
timestamp 1626908933
transform 1 0 9264 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3624
timestamp 1626908933
transform 1 0 9552 0 1 30895
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1689
timestamp 1626908933
transform 1 0 9552 0 1 30895
box -29 -23 29 23
use M1M2_PR  M1M2_PR_3564
timestamp 1626908933
transform 1 0 9552 0 1 30895
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1597
timestamp 1626908933
transform 1 0 9552 0 1 30895
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2980
timestamp 1626908933
transform 1 0 9456 0 1 30969
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1045
timestamp 1626908933
transform 1 0 9456 0 1 30969
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_25
timestamp 1626908933
transform 1 0 9984 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_382
timestamp 1626908933
transform 1 0 9984 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_29
timestamp 1626908933
transform 1 0 9888 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1020
timestamp 1626908933
transform 1 0 9888 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_500
timestamp 1626908933
transform 1 0 9984 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1222
timestamp 1626908933
transform 1 0 9984 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_431
timestamp 1626908933
transform 1 0 9600 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1029
timestamp 1626908933
transform 1 0 9600 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_37
timestamp 1626908933
transform -1 0 9600 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_99
timestamp 1626908933
transform -1 0 9600 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_216
timestamp 1626908933
transform 1 0 10100 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_864
timestamp 1626908933
transform 1 0 10100 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_216
timestamp 1626908933
transform 1 0 10100 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_864
timestamp 1626908933
transform 1 0 10100 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_132
timestamp 1626908933
transform -1 0 11232 0 -1 31968
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_63
timestamp 1626908933
transform -1 0 11232 0 -1 31968
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_501
timestamp 1626908933
transform 1 0 10464 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1223
timestamp 1626908933
transform 1 0 10464 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_411
timestamp 1626908933
transform 1 0 10080 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1009
timestamp 1626908933
transform 1 0 10080 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1177
timestamp 1626908933
transform 1 0 11300 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_529
timestamp 1626908933
transform 1 0 11300 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1177
timestamp 1626908933
transform 1 0 11300 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_529
timestamp 1626908933
transform 1 0 11300 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1042
timestamp 1626908933
transform 1 0 11232 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1019
timestamp 1626908933
transform 1 0 11232 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_51
timestamp 1626908933
transform 1 0 11232 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_28
timestamp 1626908933
transform 1 0 11232 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_986
timestamp 1626908933
transform 1 0 11328 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_985
timestamp 1626908933
transform 1 0 11328 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_388
timestamp 1626908933
transform 1 0 11328 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_387
timestamp 1626908933
transform 1 0 11328 0 -1 31968
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_192
timestamp 1626908933
transform 1 0 12500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_840
timestamp 1626908933
transform 1 0 12500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_192
timestamp 1626908933
transform 1 0 12500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_840
timestamp 1626908933
transform 1 0 12500 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_474
timestamp 1626908933
transform 1 0 11712 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_475
timestamp 1626908933
transform 1 0 11712 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1196
timestamp 1626908933
transform 1 0 11712 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1197
timestamp 1626908933
transform 1 0 11712 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_18
timestamp 1626908933
transform 1 0 12480 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_375
timestamp 1626908933
transform 1 0 12480 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_369
timestamp 1626908933
transform 1 0 12480 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_967
timestamp 1626908933
transform 1 0 12480 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_50
timestamp 1626908933
transform 1 0 12864 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1041
timestamp 1626908933
transform 1 0 12864 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_343
timestamp 1626908933
transform 1 0 13824 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_941
timestamp 1626908933
transform 1 0 13824 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_49
timestamp 1626908933
transform 1 0 13728 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1040
timestamp 1626908933
transform 1 0 13728 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_505
timestamp 1626908933
transform 1 0 13700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1153
timestamp 1626908933
transform 1 0 13700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_505
timestamp 1626908933
transform 1 0 13700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1153
timestamp 1626908933
transform 1 0 13700 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_451
timestamp 1626908933
transform 1 0 12960 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1173
timestamp 1626908933
transform 1 0 12960 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_91
timestamp 1626908933
transform 1 0 12576 0 -1 31968
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_45
timestamp 1626908933
transform 1 0 12576 0 -1 31968
box -38 -49 2726 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1146
timestamp 1626908933
transform 1 0 14208 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_424
timestamp 1626908933
transform 1 0 14208 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_24
timestamp 1626908933
transform 1 0 14976 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_381
timestamp 1626908933
transform 1 0 14976 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_168
timestamp 1626908933
transform 1 0 14900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_816
timestamp 1626908933
transform 1 0 14900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_168
timestamp 1626908933
transform 1 0 14900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_816
timestamp 1626908933
transform 1 0 14900 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_21
timestamp 1626908933
transform 1 0 15264 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_622
timestamp 1626908933
transform 1 0 15264 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_27
timestamp 1626908933
transform 1 0 15456 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_48
timestamp 1626908933
transform 1 0 15456 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1018
timestamp 1626908933
transform 1 0 15456 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1039
timestamp 1626908933
transform 1 0 15456 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_310
timestamp 1626908933
transform 1 0 15072 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_908
timestamp 1626908933
transform 1 0 15072 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_47
timestamp 1626908933
transform 1 0 16320 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1038
timestamp 1626908933
transform 1 0 16320 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_481
timestamp 1626908933
transform 1 0 16100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1129
timestamp 1626908933
transform 1 0 16100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_481
timestamp 1626908933
transform 1 0 16100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1129
timestamp 1626908933
transform 1 0 16100 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_397
timestamp 1626908933
transform 1 0 15552 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_398
timestamp 1626908933
transform 1 0 15552 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1119
timestamp 1626908933
transform 1 0 15552 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1120
timestamp 1626908933
transform 1 0 15552 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_291
timestamp 1626908933
transform 1 0 16320 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_889
timestamp 1626908933
transform 1 0 16320 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_890
timestamp 1626908933
transform 1 0 16416 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_292
timestamp 1626908933
transform 1 0 16416 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_792
timestamp 1626908933
transform 1 0 17300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_144
timestamp 1626908933
transform 1 0 17300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_792
timestamp 1626908933
transform 1 0 17300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_144
timestamp 1626908933
transform 1 0 17300 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1094
timestamp 1626908933
transform 1 0 16800 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1093
timestamp 1626908933
transform 1 0 16704 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_372
timestamp 1626908933
transform 1 0 16800 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_371
timestamp 1626908933
transform 1 0 16704 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_17
timestamp 1626908933
transform 1 0 17472 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_374
timestamp 1626908933
transform 1 0 17472 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_26
timestamp 1626908933
transform 1 0 17568 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_46
timestamp 1626908933
transform 1 0 17568 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1017
timestamp 1626908933
transform 1 0 17568 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1037
timestamp 1626908933
transform 1 0 17568 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_25
timestamp 1626908933
transform 1 0 18048 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_45
timestamp 1626908933
transform 1 0 18048 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1016
timestamp 1626908933
transform 1 0 18048 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1036
timestamp 1626908933
transform 1 0 18048 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_342
timestamp 1626908933
transform 1 0 18144 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_343
timestamp 1626908933
transform 1 0 18144 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1064
timestamp 1626908933
transform 1 0 18144 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1065
timestamp 1626908933
transform 1 0 18144 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_253
timestamp 1626908933
transform 1 0 17664 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_254
timestamp 1626908933
transform 1 0 17664 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_851
timestamp 1626908933
transform 1 0 17664 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_852
timestamp 1626908933
transform 1 0 17664 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_457
timestamp 1626908933
transform 1 0 18500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1105
timestamp 1626908933
transform 1 0 18500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_457
timestamp 1626908933
transform 1 0 18500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1105
timestamp 1626908933
transform 1 0 18500 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_30
timestamp 1626908933
transform 1 0 18912 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_631
timestamp 1626908933
transform 1 0 18912 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_24
timestamp 1626908933
transform 1 0 18912 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_44
timestamp 1626908933
transform 1 0 19104 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1015
timestamp 1626908933
transform 1 0 18912 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1035
timestamp 1626908933
transform 1 0 19104 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_233
timestamp 1626908933
transform 1 0 19008 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_831
timestamp 1626908933
transform 1 0 19008 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1038
timestamp 1626908933
transform 1 0 19200 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_316
timestamp 1626908933
transform 1 0 19200 0 1 30636
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_120
timestamp 1626908933
transform 1 0 19700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_768
timestamp 1626908933
transform 1 0 19700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_120
timestamp 1626908933
transform 1 0 19700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_768
timestamp 1626908933
transform 1 0 19700 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_23
timestamp 1626908933
transform 1 0 19968 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_380
timestamp 1626908933
transform 1 0 19968 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_23
timestamp 1626908933
transform 1 0 20160 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1014
timestamp 1626908933
transform 1 0 20160 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_303
timestamp 1626908933
transform 1 0 20064 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_315
timestamp 1626908933
transform 1 0 19392 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1025
timestamp 1626908933
transform 1 0 20064 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1037
timestamp 1626908933
transform 1 0 19392 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_43
timestamp 1626908933
transform 1 0 20832 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1034
timestamp 1626908933
transform 1 0 20832 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_433
timestamp 1626908933
transform 1 0 20900 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1081
timestamp 1626908933
transform 1 0 20900 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_433
timestamp 1626908933
transform 1 0 20900 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1081
timestamp 1626908933
transform 1 0 20900 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_292
timestamp 1626908933
transform 1 0 20640 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1014
timestamp 1626908933
transform 1 0 20640 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_199
timestamp 1626908933
transform 1 0 20928 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_209
timestamp 1626908933
transform 1 0 20256 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_797
timestamp 1626908933
transform 1 0 20928 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_807
timestamp 1626908933
transform 1 0 20256 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_20
timestamp 1626908933
transform 1 0 21408 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_621
timestamp 1626908933
transform 1 0 21408 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_22
timestamp 1626908933
transform 1 0 21600 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1013
timestamp 1626908933
transform 1 0 21600 0 -1 31968
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1835
timestamp 1626908933
transform 1 0 21840 0 1 31043
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3802
timestamp 1626908933
transform 1 0 21840 0 1 31043
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_263
timestamp 1626908933
transform 1 0 21696 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_276
timestamp 1626908933
transform 1 0 21312 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_985
timestamp 1626908933
transform 1 0 21696 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_998
timestamp 1626908933
transform 1 0 21312 0 1 30636
box -38 -49 806 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_744
timestamp 1626908933
transform 1 0 22100 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_96
timestamp 1626908933
transform 1 0 22100 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_744
timestamp 1626908933
transform 1 0 22100 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_96
timestamp 1626908933
transform 1 0 22100 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_776
timestamp 1626908933
transform 1 0 22080 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_178
timestamp 1626908933
transform 1 0 22080 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1033
timestamp 1626908933
transform 1 0 22464 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_42
timestamp 1626908933
transform 1 0 22464 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_960
timestamp 1626908933
transform 1 0 22560 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_959
timestamp 1626908933
transform 1 0 22560 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_238
timestamp 1626908933
transform 1 0 22560 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_237
timestamp 1626908933
transform 1 0 22560 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_373
timestamp 1626908933
transform 1 0 22464 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_16
timestamp 1626908933
transform 1 0 22464 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_19
timestamp 1626908933
transform 1 0 23328 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_29
timestamp 1626908933
transform 1 0 23328 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_620
timestamp 1626908933
transform 1 0 23328 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_630
timestamp 1626908933
transform 1 0 23328 0 1 30636
box -38 -49 230 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_409
timestamp 1626908933
transform 1 0 23300 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1057
timestamp 1626908933
transform 1 0 23300 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_409
timestamp 1626908933
transform 1 0 23300 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1057
timestamp 1626908933
transform 1 0 23300 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_148
timestamp 1626908933
transform 1 0 23520 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_149
timestamp 1626908933
transform 1 0 23520 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_746
timestamp 1626908933
transform 1 0 23520 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_747
timestamp 1626908933
transform 1 0 23520 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_720
timestamp 1626908933
transform 1 0 24500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_72
timestamp 1626908933
transform 1 0 24500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_720
timestamp 1626908933
transform 1 0 24500 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_72
timestamp 1626908933
transform 1 0 24500 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_929
timestamp 1626908933
transform 1 0 23904 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_928
timestamp 1626908933
transform 1 0 23904 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_207
timestamp 1626908933
transform 1 0 23904 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_206
timestamp 1626908933
transform 1 0 23904 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1966
timestamp 1626908933
transform 1 0 24864 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1012
timestamp 1626908933
transform 1 0 24672 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_975
timestamp 1626908933
transform 1 0 24864 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_21
timestamp 1626908933
transform 1 0 24672 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1197
timestamp 1626908933
transform 1 0 24672 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_596
timestamp 1626908933
transform 1 0 24672 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_724
timestamp 1626908933
transform 1 0 24768 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_126
timestamp 1626908933
transform 1 0 24768 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_22
timestamp 1626908933
transform 1 0 24960 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_379
timestamp 1626908933
transform 1 0 24960 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_41
timestamp 1626908933
transform 1 0 25056 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1032
timestamp 1626908933
transform 1 0 25056 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_385
timestamp 1626908933
transform 1 0 25700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1033
timestamp 1626908933
transform 1 0 25700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_385
timestamp 1626908933
transform 1 0 25700 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1033
timestamp 1626908933
transform 1 0 25700 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_172
timestamp 1626908933
transform 1 0 25152 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_173
timestamp 1626908933
transform 1 0 25152 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_894
timestamp 1626908933
transform 1 0 25152 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_895
timestamp 1626908933
transform 1 0 25152 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_18
timestamp 1626908933
transform 1 0 25920 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_28
timestamp 1626908933
transform 1 0 25920 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_619
timestamp 1626908933
transform 1 0 25920 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_629
timestamp 1626908933
transform 1 0 25920 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_144
timestamp 1626908933
transform 1 0 26496 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_145
timestamp 1626908933
transform 1 0 26496 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_866
timestamp 1626908933
transform 1 0 26496 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_867
timestamp 1626908933
transform 1 0 26496 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_96
timestamp 1626908933
transform 1 0 26112 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_97
timestamp 1626908933
transform 1 0 26112 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_694
timestamp 1626908933
transform 1 0 26112 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_695
timestamp 1626908933
transform 1 0 26112 0 1 30636
box -38 -49 422 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_48
timestamp 1626908933
transform 1 0 26900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_696
timestamp 1626908933
transform 1 0 26900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_48
timestamp 1626908933
transform 1 0 26900 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_696
timestamp 1626908933
transform 1 0 26900 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_20
timestamp 1626908933
transform 1 0 27264 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_40
timestamp 1626908933
transform 1 0 27264 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_978
timestamp 1626908933
transform 1 0 27360 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1011
timestamp 1626908933
transform 1 0 27264 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1031
timestamp 1626908933
transform 1 0 27264 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1969
timestamp 1626908933
transform 1 0 27360 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_79
timestamp 1626908933
transform 1 0 27360 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_677
timestamp 1626908933
transform 1 0 27360 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_618
timestamp 1626908933
transform 1 0 27552 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_17
timestamp 1626908933
transform 1 0 27552 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_372
timestamp 1626908933
transform 1 0 27456 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_15
timestamp 1626908933
transform 1 0 27456 0 -1 31968
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1009
timestamp 1626908933
transform 1 0 28100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_361
timestamp 1626908933
transform 1 0 28100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1009
timestamp 1626908933
transform 1 0 28100 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_361
timestamp 1626908933
transform 1 0 28100 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_834
timestamp 1626908933
transform 1 0 27744 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_833
timestamp 1626908933
transform 1 0 27744 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_112
timestamp 1626908933
transform 1 0 27744 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_111
timestamp 1626908933
transform 1 0 27744 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_19
timestamp 1626908933
transform 1 0 28896 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_39
timestamp 1626908933
transform 1 0 28896 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1010
timestamp 1626908933
transform 1 0 28896 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1030
timestamp 1626908933
transform 1 0 28896 0 1 30636
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_24
timestamp 1626908933
transform 1 0 29300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_672
timestamp 1626908933
transform 1 0 29300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_24
timestamp 1626908933
transform 1 0 29300 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_672
timestamp 1626908933
transform 1 0 29300 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_77
timestamp 1626908933
transform 1 0 28992 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_78
timestamp 1626908933
transform 1 0 28992 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_799
timestamp 1626908933
transform 1 0 28992 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_800
timestamp 1626908933
transform 1 0 28992 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_51
timestamp 1626908933
transform 1 0 28512 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_52
timestamp 1626908933
transform 1 0 28512 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_649
timestamp 1626908933
transform 1 0 28512 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_650
timestamp 1626908933
transform 1 0 28512 0 1 30636
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_16
timestamp 1626908933
transform 1 0 29760 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_617
timestamp 1626908933
transform 1 0 29760 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_38
timestamp 1626908933
transform 1 0 29760 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1029
timestamp 1626908933
transform 1 0 29760 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_21
timestamp 1626908933
transform 1 0 29952 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_378
timestamp 1626908933
transform 1 0 29952 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_27
timestamp 1626908933
transform 1 0 30048 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_628
timestamp 1626908933
transform 1 0 30048 0 1 30636
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_976
timestamp 1626908933
transform 1 0 29856 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1967
timestamp 1626908933
transform 1 0 29856 0 1 30636
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1829
timestamp 1626908933
transform 1 0 30096 0 1 31191
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3796
timestamp 1626908933
transform 1 0 30096 0 1 31191
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_23
timestamp 1626908933
transform 1 0 29952 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_621
timestamp 1626908933
transform 1 0 29952 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1028
timestamp 1626908933
transform 1 0 30240 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_37
timestamp 1626908933
transform 1 0 30240 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_753
timestamp 1626908933
transform 1 0 30336 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_752
timestamp 1626908933
transform 1 0 30336 0 -1 31968
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_31
timestamp 1626908933
transform 1 0 30336 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_30
timestamp 1626908933
transform 1 0 30336 0 -1 31968
box -38 -49 806 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_337
timestamp 1626908933
transform 1 0 30500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_985
timestamp 1626908933
transform 1 0 30500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_337
timestamp 1626908933
transform 1 0 30500 0 1 30636
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_985
timestamp 1626908933
transform 1 0 30500 0 1 30636
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_36
timestamp 1626908933
transform 1 0 31104 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1027
timestamp 1626908933
transform 1 0 31104 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_0
timestamp 1626908933
transform 1 0 31200 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_722
timestamp 1626908933
transform 1 0 31200 0 1 30636
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1
timestamp 1626908933
transform 1 0 31104 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_599
timestamp 1626908933
transform 1 0 31104 0 -1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_18
timestamp 1626908933
transform 1 0 31488 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1009
timestamp 1626908933
transform 1 0 31488 0 -1 31968
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_648
timestamp 1626908933
transform 1 0 31700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_0
timestamp 1626908933
transform 1 0 31700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_648
timestamp 1626908933
transform 1 0 31700 0 1 31302
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_0
timestamp 1626908933
transform 1 0 31700 0 1 31302
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1970
timestamp 1626908933
transform 1 0 31584 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_979
timestamp 1626908933
transform 1 0 31584 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1199
timestamp 1626908933
transform 1 0 31776 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_598
timestamp 1626908933
transform 1 0 31776 0 -1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_371
timestamp 1626908933
transform 1 0 31680 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_14
timestamp 1626908933
transform 1 0 31680 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_977
timestamp 1626908933
transform 1 0 31968 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_980
timestamp 1626908933
transform 1 0 31968 0 -1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1968
timestamp 1626908933
transform 1 0 31968 0 1 30636
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1971
timestamp 1626908933
transform 1 0 31968 0 -1 31968
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1828
timestamp 1626908933
transform 1 0 32016 0 1 31191
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3795
timestamp 1626908933
transform 1 0 32016 0 1 31191
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1972
timestamp 1626908933
transform 1 0 192 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1008
timestamp 1626908933
transform 1 0 384 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_981
timestamp 1626908933
transform 1 0 192 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_17
timestamp 1626908933
transform 1 0 384 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1200
timestamp 1626908933
transform 1 0 0 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_599
timestamp 1626908933
transform 1 0 0 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_370
timestamp 1626908933
transform 1 0 288 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_13
timestamp 1626908933
transform 1 0 288 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1184
timestamp 1626908933
transform 1 0 480 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1183
timestamp 1626908933
transform 1 0 864 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_586
timestamp 1626908933
transform 1 0 480 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_585
timestamp 1626908933
transform 1 0 864 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1159
timestamp 1626908933
transform 1 0 1248 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_561
timestamp 1626908933
transform 1 0 1248 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1272
timestamp 1626908933
transform 1 0 1700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_624
timestamp 1626908933
transform 1 0 1700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1272
timestamp 1626908933
transform 1 0 1700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_624
timestamp 1626908933
transform 1 0 1700 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1154
timestamp 1626908933
transform 1 0 1632 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_556
timestamp 1626908933
transform 1 0 1632 0 1 31968
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2172
timestamp 1626908933
transform 1 0 2064 0 1 31635
box -32 -32 32 32
use M1M2_PR  M1M2_PR_205
timestamp 1626908933
transform 1 0 2064 0 1 31635
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1150
timestamp 1626908933
transform 1 0 2016 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_552
timestamp 1626908933
transform 1 0 2016 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1007
timestamp 1626908933
transform 1 0 2400 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_16
timestamp 1626908933
transform 1 0 2400 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_616
timestamp 1626908933
transform 1 0 2592 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_15
timestamp 1626908933
transform 1 0 2592 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_369
timestamp 1626908933
transform 1 0 2496 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_12
timestamp 1626908933
transform 1 0 2496 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_615
timestamp 1626908933
transform 1 0 3168 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_14
timestamp 1626908933
transform 1 0 3168 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1143
timestamp 1626908933
transform 1 0 2784 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_545
timestamp 1626908933
transform 1 0 2784 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1006
timestamp 1626908933
transform 1 0 3360 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_15
timestamp 1626908933
transform 1 0 3360 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1128
timestamp 1626908933
transform 1 0 3456 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_530
timestamp 1626908933
transform 1 0 3456 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1248
timestamp 1626908933
transform 1 0 4100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_600
timestamp 1626908933
transform 1 0 4100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1248
timestamp 1626908933
transform 1 0 4100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_600
timestamp 1626908933
transform 1 0 4100 0 1 31968
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2159
timestamp 1626908933
transform 1 0 4080 0 1 31635
box -29 -23 29 23
use L1M1_PR  L1M1_PR_224
timestamp 1626908933
transform 1 0 4080 0 1 31635
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1123
timestamp 1626908933
transform 1 0 3840 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_525
timestamp 1626908933
transform 1 0 3840 0 1 31968
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2992
timestamp 1626908933
transform 1 0 4272 0 1 31561
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1057
timestamp 1626908933
transform 1 0 4272 0 1 31561
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2171
timestamp 1626908933
transform 1 0 4176 0 1 31635
box -32 -32 32 32
use M1M2_PR  M1M2_PR_204
timestamp 1626908933
transform 1 0 4176 0 1 31635
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1121
timestamp 1626908933
transform 1 0 4224 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1111
timestamp 1626908933
transform 1 0 4608 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_523
timestamp 1626908933
transform 1 0 4224 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_513
timestamp 1626908933
transform 1 0 4608 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_368
timestamp 1626908933
transform 1 0 4992 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_11
timestamp 1626908933
transform 1 0 4992 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1005
timestamp 1626908933
transform 1 0 5280 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_14
timestamp 1626908933
transform 1 0 5280 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_614
timestamp 1626908933
transform 1 0 5088 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_13
timestamp 1626908933
transform 1 0 5088 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1097
timestamp 1626908933
transform 1 0 5376 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_499
timestamp 1626908933
transform 1 0 5376 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1095
timestamp 1626908933
transform 1 0 5760 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_497
timestamp 1626908933
transform 1 0 5760 0 1 31968
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2991
timestamp 1626908933
transform 1 0 6384 0 1 31561
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1056
timestamp 1626908933
transform 1 0 6384 0 1 31561
box -29 -23 29 23
use M1M2_PR  M1M2_PR_2964
timestamp 1626908933
transform 1 0 6288 0 1 31413
box -32 -32 32 32
use M1M2_PR  M1M2_PR_997
timestamp 1626908933
transform 1 0 6288 0 1 31413
box -32 -32 32 32
use fine_freq_track_VIA1  fine_freq_track_VIA1_1224
timestamp 1626908933
transform 1 0 6500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_576
timestamp 1626908933
transform 1 0 6500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1224
timestamp 1626908933
transform 1 0 6500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_576
timestamp 1626908933
transform 1 0 6500 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1004
timestamp 1626908933
transform 1 0 6336 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_13
timestamp 1626908933
transform 1 0 6336 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_482
timestamp 1626908933
transform 1 0 6432 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1080
timestamp 1626908933
transform 1 0 6432 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_12
timestamp 1626908933
transform 1 0 6144 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_613
timestamp 1626908933
transform 1 0 6144 0 1 31968
box -38 -49 230 715
use M1M2_PR  M1M2_PR_989
timestamp 1626908933
transform 1 0 6768 0 1 31413
box -32 -32 32 32
use M1M2_PR  M1M2_PR_993
timestamp 1626908933
transform 1 0 6576 0 1 31561
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2956
timestamp 1626908933
transform 1 0 6768 0 1 31413
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2960
timestamp 1626908933
transform 1 0 6576 0 1 31561
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1053
timestamp 1626908933
transform 1 0 6768 0 1 31413
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1058
timestamp 1626908933
transform 1 0 6576 0 1 31413
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2988
timestamp 1626908933
transform 1 0 6768 0 1 31413
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2993
timestamp 1626908933
transform 1 0 6576 0 1 31413
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_476
timestamp 1626908933
transform 1 0 6816 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1074
timestamp 1626908933
transform 1 0 6816 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_612
timestamp 1626908933
transform 1 0 7200 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_11
timestamp 1626908933
transform 1 0 7200 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1973
timestamp 1626908933
transform 1 0 7392 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_982
timestamp 1626908933
transform 1 0 7392 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1057
timestamp 1626908933
transform 1 0 7584 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_459
timestamp 1626908933
transform 1 0 7584 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_367
timestamp 1626908933
transform 1 0 7488 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_10
timestamp 1626908933
transform 1 0 7488 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1054
timestamp 1626908933
transform 1 0 7968 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_456
timestamp 1626908933
transform 1 0 7968 0 1 31968
box -38 -49 422 715
use M1M2_PR  M1M2_PR_982
timestamp 1626908933
transform 1 0 8688 0 1 31635
box -32 -32 32 32
use M1M2_PR  M1M2_PR_986
timestamp 1626908933
transform 1 0 8304 0 1 31413
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2949
timestamp 1626908933
transform 1 0 8688 0 1 31635
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2953
timestamp 1626908933
transform 1 0 8304 0 1 31413
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1046
timestamp 1626908933
transform 1 0 8592 0 1 31635
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1048
timestamp 1626908933
transform 1 0 8688 0 1 31413
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2981
timestamp 1626908933
transform 1 0 8592 0 1 31635
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2983
timestamp 1626908933
transform 1 0 8688 0 1 31413
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_442
timestamp 1626908933
transform 1 0 8736 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_453
timestamp 1626908933
transform 1 0 8352 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1040
timestamp 1626908933
transform 1 0 8736 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1051
timestamp 1626908933
transform 1 0 8352 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1200
timestamp 1626908933
transform 1 0 8900 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_552
timestamp 1626908933
transform 1 0 8900 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1200
timestamp 1626908933
transform 1 0 8900 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_552
timestamp 1626908933
transform 1 0 8900 0 1 31968
box -100 -49 100 49
use L1M1_PR  L1M1_PR_3625
timestamp 1626908933
transform 1 0 8784 0 1 31635
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1690
timestamp 1626908933
transform 1 0 8784 0 1 31635
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1038
timestamp 1626908933
transform 1 0 9120 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_440
timestamp 1626908933
transform 1 0 9120 0 1 31968
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3563
timestamp 1626908933
transform 1 0 9552 0 1 31635
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1596
timestamp 1626908933
transform 1 0 9552 0 1 31635
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1003
timestamp 1626908933
transform 1 0 9504 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_12
timestamp 1626908933
transform 1 0 9504 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1028
timestamp 1626908933
transform 1 0 9600 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_430
timestamp 1626908933
transform 1 0 9600 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1002
timestamp 1626908933
transform 1 0 10080 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_11
timestamp 1626908933
transform 1 0 10080 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_366
timestamp 1626908933
transform 1 0 9984 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_9
timestamp 1626908933
transform 1 0 9984 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1008
timestamp 1626908933
transform 1 0 10176 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1005
timestamp 1626908933
transform 1 0 10560 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_410
timestamp 1626908933
transform 1 0 10176 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_407
timestamp 1626908933
transform 1 0 10560 0 1 31968
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3623
timestamp 1626908933
transform 1 0 10704 0 1 31635
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1688
timestamp 1626908933
transform 1 0 10704 0 1 31635
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1002
timestamp 1626908933
transform 1 0 10944 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_404
timestamp 1626908933
transform 1 0 10944 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1176
timestamp 1626908933
transform 1 0 11300 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_528
timestamp 1626908933
transform 1 0 11300 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1176
timestamp 1626908933
transform 1 0 11300 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_528
timestamp 1626908933
transform 1 0 11300 0 1 31968
box -100 -49 100 49
use L1M1_PR  L1M1_PR_2150
timestamp 1626908933
transform 1 0 11280 0 1 31487
box -29 -23 29 23
use L1M1_PR  L1M1_PR_215
timestamp 1626908933
transform 1 0 11280 0 1 31487
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_984
timestamp 1626908933
transform 1 0 11328 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_386
timestamp 1626908933
transform 1 0 11328 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_982
timestamp 1626908933
transform 1 0 11712 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_384
timestamp 1626908933
transform 1 0 11712 0 1 31968
box -38 -49 422 715
use M1M2_PR  M1M2_PR_3587
timestamp 1626908933
transform 1 0 12336 0 1 31635
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1620
timestamp 1626908933
transform 1 0 12336 0 1 31635
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_973
timestamp 1626908933
transform 1 0 12096 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_375
timestamp 1626908933
transform 1 0 12096 0 1 31968
box -38 -49 422 715
use L1M1_PR  L1M1_PR_3622
timestamp 1626908933
transform 1 0 12624 0 1 31709
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1687
timestamp 1626908933
transform 1 0 12624 0 1 31709
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_611
timestamp 1626908933
transform 1 0 12576 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_10
timestamp 1626908933
transform 1 0 12576 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_953
timestamp 1626908933
transform 1 0 12768 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_355
timestamp 1626908933
transform 1 0 12768 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_365
timestamp 1626908933
transform 1 0 12480 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_8
timestamp 1626908933
transform 1 0 12480 0 1 31968
box -38 -49 134 715
use L1M1_PR  L1M1_PR_3641
timestamp 1626908933
transform 1 0 13008 0 1 31635
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1706
timestamp 1626908933
transform 1 0 13008 0 1 31635
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_948
timestamp 1626908933
transform 1 0 13152 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_350
timestamp 1626908933
transform 1 0 13152 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1152
timestamp 1626908933
transform 1 0 13700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_504
timestamp 1626908933
transform 1 0 13700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1152
timestamp 1626908933
transform 1 0 13700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_504
timestamp 1626908933
transform 1 0 13700 0 1 31968
box -100 -49 100 49
use M1M2_PR  M1M2_PR_3683
timestamp 1626908933
transform 1 0 13488 0 1 31561
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1716
timestamp 1626908933
transform 1 0 13488 0 1 31561
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_946
timestamp 1626908933
transform 1 0 13536 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_348
timestamp 1626908933
transform 1 0 13536 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_940
timestamp 1626908933
transform 1 0 13920 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_342
timestamp 1626908933
transform 1 0 13920 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_610
timestamp 1626908933
transform 1 0 14688 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_9
timestamp 1626908933
transform 1 0 14688 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_937
timestamp 1626908933
transform 1 0 14304 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_339
timestamp 1626908933
transform 1 0 14304 0 1 31968
box -38 -49 422 715
use L1M1_PR  L1M1_PR_2149
timestamp 1626908933
transform 1 0 14832 0 1 31487
box -29 -23 29 23
use L1M1_PR  L1M1_PR_214
timestamp 1626908933
transform 1 0 14832 0 1 31487
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1974
timestamp 1626908933
transform 1 0 14880 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_983
timestamp 1626908933
transform 1 0 14880 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_907
timestamp 1626908933
transform 1 0 15072 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_309
timestamp 1626908933
transform 1 0 15072 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_364
timestamp 1626908933
transform 1 0 14976 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_7
timestamp 1626908933
transform 1 0 14976 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_906
timestamp 1626908933
transform 1 0 15456 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_308
timestamp 1626908933
transform 1 0 15456 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_10
timestamp 1626908933
transform 1 0 16032 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1001
timestamp 1626908933
transform 1 0 16032 0 1 31968
box -38 -49 134 715
use fine_freq_track_VIA0  fine_freq_track_VIA0_480
timestamp 1626908933
transform 1 0 16100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1128
timestamp 1626908933
transform 1 0 16100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_480
timestamp 1626908933
transform 1 0 16100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_1128
timestamp 1626908933
transform 1 0 16100 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_300
timestamp 1626908933
transform 1 0 16128 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_898
timestamp 1626908933
transform 1 0 16128 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_8
timestamp 1626908933
transform 1 0 15840 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_609
timestamp 1626908933
transform 1 0 15840 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_888
timestamp 1626908933
transform 1 0 16512 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_290
timestamp 1626908933
transform 1 0 16512 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_883
timestamp 1626908933
transform 1 0 16896 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_285
timestamp 1626908933
transform 1 0 16896 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1975
timestamp 1626908933
transform 1 0 17376 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1000
timestamp 1626908933
transform 1 0 17280 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_984
timestamp 1626908933
transform 1 0 17376 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_9
timestamp 1626908933
transform 1 0 17280 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_363
timestamp 1626908933
transform 1 0 17472 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_6
timestamp 1626908933
transform 1 0 17472 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_999
timestamp 1626908933
transform 1 0 17568 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_8
timestamp 1626908933
transform 1 0 17568 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_850
timestamp 1626908933
transform 1 0 17664 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_252
timestamp 1626908933
transform 1 0 17664 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_848
timestamp 1626908933
transform 1 0 18048 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_845
timestamp 1626908933
transform 1 0 18432 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_250
timestamp 1626908933
transform 1 0 18048 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_247
timestamp 1626908933
transform 1 0 18432 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1104
timestamp 1626908933
transform 1 0 18500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_456
timestamp 1626908933
transform 1 0 18500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1104
timestamp 1626908933
transform 1 0 18500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_456
timestamp 1626908933
transform 1 0 18500 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_841
timestamp 1626908933
transform 1 0 18816 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_243
timestamp 1626908933
transform 1 0 18816 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_608
timestamp 1626908933
transform 1 0 19200 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_7
timestamp 1626908933
transform 1 0 19200 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_998
timestamp 1626908933
transform 1 0 19392 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_7
timestamp 1626908933
transform 1 0 19392 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_823
timestamp 1626908933
transform 1 0 19488 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_225
timestamp 1626908933
transform 1 0 19488 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1976
timestamp 1626908933
transform 1 0 19872 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_985
timestamp 1626908933
transform 1 0 19872 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_607
timestamp 1626908933
transform 1 0 20064 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_6
timestamp 1626908933
transform 1 0 20064 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_806
timestamp 1626908933
transform 1 0 20256 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_208
timestamp 1626908933
transform 1 0 20256 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_362
timestamp 1626908933
transform 1 0 19968 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_5
timestamp 1626908933
transform 1 0 19968 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_805
timestamp 1626908933
transform 1 0 20640 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_207
timestamp 1626908933
transform 1 0 20640 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1080
timestamp 1626908933
transform 1 0 20900 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_432
timestamp 1626908933
transform 1 0 20900 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1080
timestamp 1626908933
transform 1 0 20900 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_432
timestamp 1626908933
transform 1 0 20900 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_796
timestamp 1626908933
transform 1 0 21024 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_198
timestamp 1626908933
transform 1 0 21024 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_792
timestamp 1626908933
transform 1 0 21408 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_194
timestamp 1626908933
transform 1 0 21408 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_790
timestamp 1626908933
transform 1 0 21792 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_192
timestamp 1626908933
transform 1 0 21792 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1977
timestamp 1626908933
transform 1 0 22368 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_986
timestamp 1626908933
transform 1 0 22368 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_606
timestamp 1626908933
transform 1 0 22176 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_605
timestamp 1626908933
transform 1 0 22560 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_5
timestamp 1626908933
transform 1 0 22176 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_4
timestamp 1626908933
transform 1 0 22560 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_361
timestamp 1626908933
transform 1 0 22464 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_4
timestamp 1626908933
transform 1 0 22464 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_997
timestamp 1626908933
transform 1 0 22752 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_6
timestamp 1626908933
transform 1 0 22752 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_765
timestamp 1626908933
transform 1 0 22848 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_167
timestamp 1626908933
transform 1 0 22848 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1056
timestamp 1626908933
transform 1 0 23300 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_408
timestamp 1626908933
transform 1 0 23300 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1056
timestamp 1626908933
transform 1 0 23300 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_408
timestamp 1626908933
transform 1 0 23300 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_764
timestamp 1626908933
transform 1 0 23232 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_166
timestamp 1626908933
transform 1 0 23232 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_745
timestamp 1626908933
transform 1 0 23616 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_147
timestamp 1626908933
transform 1 0 23616 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_743
timestamp 1626908933
transform 1 0 24000 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_739
timestamp 1626908933
transform 1 0 24384 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_145
timestamp 1626908933
transform 1 0 24000 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_141
timestamp 1626908933
transform 1 0 24384 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1978
timestamp 1626908933
transform 1 0 24864 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_996
timestamp 1626908933
transform 1 0 24768 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_987
timestamp 1626908933
transform 1 0 24864 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_5
timestamp 1626908933
transform 1 0 24768 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_995
timestamp 1626908933
transform 1 0 25056 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_4
timestamp 1626908933
transform 1 0 25056 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_718
timestamp 1626908933
transform 1 0 25152 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_120
timestamp 1626908933
transform 1 0 25152 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_360
timestamp 1626908933
transform 1 0 24960 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1626908933
transform 1 0 24960 0 1 31968
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1032
timestamp 1626908933
transform 1 0 25700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_384
timestamp 1626908933
transform 1 0 25700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1032
timestamp 1626908933
transform 1 0 25700 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_384
timestamp 1626908933
transform 1 0 25700 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_994
timestamp 1626908933
transform 1 0 25728 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_3
timestamp 1626908933
transform 1 0 25728 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_604
timestamp 1626908933
transform 1 0 25536 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_3
timestamp 1626908933
transform 1 0 25536 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_714
timestamp 1626908933
transform 1 0 25824 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_693
timestamp 1626908933
transform 1 0 26208 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_116
timestamp 1626908933
transform 1 0 25824 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_95
timestamp 1626908933
transform 1 0 26208 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_691
timestamp 1626908933
transform 1 0 26592 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_93
timestamp 1626908933
transform 1 0 26592 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_688
timestamp 1626908933
transform 1 0 26976 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_90
timestamp 1626908933
transform 1 0 26976 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1979
timestamp 1626908933
transform 1 0 27360 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_988
timestamp 1626908933
transform 1 0 27360 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_603
timestamp 1626908933
transform 1 0 27552 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_2
timestamp 1626908933
transform 1 0 27552 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_359
timestamp 1626908933
transform 1 0 27456 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1626908933
transform 1 0 27456 0 1 31968
box -38 -49 134 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_1008
timestamp 1626908933
transform 1 0 28100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_360
timestamp 1626908933
transform 1 0 28100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_1008
timestamp 1626908933
transform 1 0 28100 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_360
timestamp 1626908933
transform 1 0 28100 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_674
timestamp 1626908933
transform 1 0 27744 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_76
timestamp 1626908933
transform 1 0 27744 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_670
timestamp 1626908933
transform 1 0 28128 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_648
timestamp 1626908933
transform 1 0 28512 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_72
timestamp 1626908933
transform 1 0 28128 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_50
timestamp 1626908933
transform 1 0 28512 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_602
timestamp 1626908933
transform 1 0 28896 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1
timestamp 1626908933
transform 1 0 28896 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_993
timestamp 1626908933
transform 1 0 29088 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_2
timestamp 1626908933
transform 1 0 29088 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_644
timestamp 1626908933
transform 1 0 29184 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_46
timestamp 1626908933
transform 1 0 29184 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_637
timestamp 1626908933
transform 1 0 29568 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_39
timestamp 1626908933
transform 1 0 29568 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_358
timestamp 1626908933
transform 1 0 29952 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1626908933
transform 1 0 29952 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_992
timestamp 1626908933
transform 1 0 30240 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1
timestamp 1626908933
transform 1 0 30240 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_601
timestamp 1626908933
transform 1 0 30048 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_0
timestamp 1626908933
transform 1 0 30048 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_620
timestamp 1626908933
transform 1 0 30336 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_22
timestamp 1626908933
transform 1 0 30336 0 1 31968
box -38 -49 422 715
use fine_freq_track_VIA1  fine_freq_track_VIA1_984
timestamp 1626908933
transform 1 0 30500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA1  fine_freq_track_VIA1_336
timestamp 1626908933
transform 1 0 30500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_984
timestamp 1626908933
transform 1 0 30500 0 1 31968
box -100 -49 100 49
use fine_freq_track_VIA0  fine_freq_track_VIA0_336
timestamp 1626908933
transform 1 0 30500 0 1 31968
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_616
timestamp 1626908933
transform 1 0 30720 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_18
timestamp 1626908933
transform 1 0 30720 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_598
timestamp 1626908933
transform 1 0 31104 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_0
timestamp 1626908933
transform 1 0 31104 0 1 31968
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1980
timestamp 1626908933
transform 1 0 31584 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_991
timestamp 1626908933
transform 1 0 31488 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_989
timestamp 1626908933
transform 1 0 31584 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_0
timestamp 1626908933
transform 1 0 31488 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1201
timestamp 1626908933
transform 1 0 31776 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_600
timestamp 1626908933
transform 1 0 31776 0 1 31968
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_357
timestamp 1626908933
transform 1 0 31680 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0
timestamp 1626908933
transform 1 0 31680 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1981
timestamp 1626908933
transform 1 0 31968 0 1 31968
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_990
timestamp 1626908933
transform 1 0 31968 0 1 31968
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1833
timestamp 1626908933
transform 1 0 48 0 1 32375
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3800
timestamp 1626908933
transform 1 0 48 0 1 32375
box -32 -32 32 32
use fine_freq_track_VIA2  fine_freq_track_VIA2_13
timestamp 1626908933
transform 1 0 500 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_40
timestamp 1626908933
transform 1 0 500 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_13
timestamp 1626908933
transform 1 0 500 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_40
timestamp 1626908933
transform 1 0 500 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_11
timestamp 1626908933
transform 1 0 5300 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_12
timestamp 1626908933
transform 1 0 2900 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_38
timestamp 1626908933
transform 1 0 5300 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_39
timestamp 1626908933
transform 1 0 2900 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_11
timestamp 1626908933
transform 1 0 5300 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_12
timestamp 1626908933
transform 1 0 2900 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_38
timestamp 1626908933
transform 1 0 5300 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_39
timestamp 1626908933
transform 1 0 2900 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_10
timestamp 1626908933
transform 1 0 7700 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_37
timestamp 1626908933
transform 1 0 7700 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_10
timestamp 1626908933
transform 1 0 7700 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_37
timestamp 1626908933
transform 1 0 7700 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_9
timestamp 1626908933
transform 1 0 10100 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_36
timestamp 1626908933
transform 1 0 10100 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_9
timestamp 1626908933
transform 1 0 10100 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_36
timestamp 1626908933
transform 1 0 10100 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_8
timestamp 1626908933
transform 1 0 12500 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_35
timestamp 1626908933
transform 1 0 12500 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_8
timestamp 1626908933
transform 1 0 12500 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_35
timestamp 1626908933
transform 1 0 12500 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_7
timestamp 1626908933
transform 1 0 14900 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_34
timestamp 1626908933
transform 1 0 14900 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_7
timestamp 1626908933
transform 1 0 14900 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_34
timestamp 1626908933
transform 1 0 14900 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_6
timestamp 1626908933
transform 1 0 17300 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_33
timestamp 1626908933
transform 1 0 17300 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_6
timestamp 1626908933
transform 1 0 17300 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_33
timestamp 1626908933
transform 1 0 17300 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_4
timestamp 1626908933
transform 1 0 22100 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_5
timestamp 1626908933
transform 1 0 19700 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_31
timestamp 1626908933
transform 1 0 22100 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_32
timestamp 1626908933
transform 1 0 19700 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_4
timestamp 1626908933
transform 1 0 22100 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_5
timestamp 1626908933
transform 1 0 19700 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_31
timestamp 1626908933
transform 1 0 22100 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_32
timestamp 1626908933
transform 1 0 19700 0 1 32611
box -100 -26 100 26
use M1M2_PR  M1M2_PR_1832
timestamp 1626908933
transform 1 0 24720 0 1 32301
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3799
timestamp 1626908933
transform 1 0 24720 0 1 32301
box -32 -32 32 32
use fine_freq_track_VIA2  fine_freq_track_VIA2_3
timestamp 1626908933
transform 1 0 24500 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_30
timestamp 1626908933
transform 1 0 24500 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_3
timestamp 1626908933
transform 1 0 24500 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_30
timestamp 1626908933
transform 1 0 24500 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_2
timestamp 1626908933
transform 1 0 26900 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_29
timestamp 1626908933
transform 1 0 26900 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_2
timestamp 1626908933
transform 1 0 26900 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_29
timestamp 1626908933
transform 1 0 26900 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_1
timestamp 1626908933
transform 1 0 29300 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_28
timestamp 1626908933
transform 1 0 29300 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_1
timestamp 1626908933
transform 1 0 29300 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_28
timestamp 1626908933
transform 1 0 29300 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA2  fine_freq_track_VIA2_0
timestamp 1626908933
transform 1 0 31700 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA2  fine_freq_track_VIA2_27
timestamp 1626908933
transform 1 0 31700 0 1 32618
box -100 -33 100 33
use fine_freq_track_VIA3  fine_freq_track_VIA3_0
timestamp 1626908933
transform 1 0 31700 0 1 32611
box -100 -26 100 26
use fine_freq_track_VIA3  fine_freq_track_VIA3_27
timestamp 1626908933
transform 1 0 31700 0 1 32611
box -100 -26 100 26
<< labels >>
rlabel metal2 s 0 17635 97 17663 4 clk_out
port 1 nsew
rlabel metal2 s 0 23 97 51 4 div_ratio_half[5]
port 2 nsew
rlabel metal2 s 0 1355 97 1383 4 div_ratio_half[4]
port 3 nsew
rlabel metal2 s 0 2687 97 2715 4 div_ratio_half[3]
port 4 nsew
rlabel metal2 s 0 4093 97 4121 4 div_ratio_half[2]
port 5 nsew
rlabel metal2 s 0 5425 97 5453 4 div_ratio_half[1]
port 6 nsew
rlabel metal2 s 0 6757 97 6785 4 div_ratio_half[0]
port 7 nsew
rlabel metal2 s 0 16303 97 16331 4 ref_clk
port 8 nsew
rlabel metal2 s 0 8089 97 8117 4 rst
port 9 nsew
rlabel metal2 s 0 9495 97 9523 4 aux_osc_en
port 10 nsew
rlabel metal2 s 0 10827 97 10855 4 fftl_en
port 11 nsew
rlabel metal2 s 0 12233 97 12261 4 fine_control_avg_window_select[4]
port 12 nsew
rlabel metal2 s 0 13565 97 13593 4 fine_control_avg_window_select[3]
port 13 nsew
rlabel metal2 s 0 18967 97 18995 4 fine_control_avg_window_select[2]
port 14 nsew
rlabel metal2 s 0 20373 97 20401 4 fine_control_avg_window_select[1]
port 15 nsew
rlabel metal2 s 0 21705 97 21733 4 fine_control_avg_window_select[0]
port 16 nsew
rlabel metal2 s 0 23037 97 23065 4 fine_con_step_size[3]
port 17 nsew
rlabel metal2 s 0 24369 97 24397 4 fine_con_step_size[2]
port 18 nsew
rlabel metal2 s 0 25775 97 25803 4 fine_con_step_size[1]
port 19 nsew
rlabel metal2 s 0 27107 97 27135 4 fine_con_step_size[0]
port 20 nsew
rlabel metal2 s 0 28439 97 28467 4 manual_control_osc[12]
port 21 nsew
rlabel metal2 s 0 29845 97 29873 4 manual_control_osc[11]
port 22 nsew
rlabel metal2 s 0 31177 97 31205 4 manual_control_osc[10]
port 23 nsew
rlabel metal2 s 0 32509 97 32537 4 manual_control_osc[9]
port 24 nsew
rlabel metal2 s 31967 32583 32064 32611 4 manual_control_osc[8]
port 25 nsew
rlabel metal2 s 31967 31103 32064 31131 4 manual_control_osc[7]
port 26 nsew
rlabel metal2 s 31967 29623 32064 29651 4 manual_control_osc[6]
port 27 nsew
rlabel metal2 s 31967 28143 32064 28171 4 manual_control_osc[5]
port 28 nsew
rlabel metal2 s 31967 26663 32064 26691 4 manual_control_osc[4]
port 29 nsew
rlabel metal2 s 31967 25183 32064 25211 4 manual_control_osc[3]
port 30 nsew
rlabel metal2 s 31967 23703 32064 23731 4 manual_control_osc[2]
port 31 nsew
rlabel metal2 s 31967 22223 32064 22251 4 manual_control_osc[1]
port 32 nsew
rlabel metal2 s 31967 20743 32064 20771 4 manual_control_osc[0]
port 33 nsew
rlabel metal2 s 0 14897 97 14925 4 aux_clk_out
port 34 nsew
rlabel metal2 s 31967 19263 32064 19291 4 out_star
port 35 nsew
rlabel metal2 s 31967 17783 32064 17811 4 osc_fine_con_final[12]
port 36 nsew
rlabel metal2 s 31967 16303 32064 16331 4 osc_fine_con_final[11]
port 37 nsew
rlabel metal2 s 31967 14823 32064 14851 4 osc_fine_con_final[10]
port 38 nsew
rlabel metal2 s 31967 13343 32064 13371 4 osc_fine_con_final[9]
port 39 nsew
rlabel metal2 s 31967 11863 32064 11891 4 osc_fine_con_final[8]
port 40 nsew
rlabel metal2 s 31967 10383 32064 10411 4 osc_fine_con_final[7]
port 41 nsew
rlabel metal2 s 31967 8903 32064 8931 4 osc_fine_con_final[6]
port 42 nsew
rlabel metal2 s 31967 7423 32064 7451 4 osc_fine_con_final[5]
port 43 nsew
rlabel metal2 s 31967 5943 32064 5971 4 osc_fine_con_final[4]
port 44 nsew
rlabel metal2 s 31967 4463 32064 4491 4 osc_fine_con_final[3]
port 45 nsew
rlabel metal2 s 31967 2983 32064 3011 4 osc_fine_con_final[2]
port 46 nsew
rlabel metal2 s 31967 1503 32064 1531 4 osc_fine_con_final[1]
port 47 nsew
rlabel metal2 s 31967 23 32064 51 4 osc_fine_con_final[0]
port 48 nsew
rlabel metal3 s 1600 0 1800 200 4 DVSS:
port 49 nsew
rlabel metal3 s 1600 32434 1800 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 4000 0 4200 200 4 DVSS:
port 49 nsew
rlabel metal3 s 4000 32434 4200 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 6400 0 6600 200 4 DVSS:
port 49 nsew
rlabel metal3 s 6400 32434 6600 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 8800 0 9000 200 4 DVSS:
port 49 nsew
rlabel metal3 s 8800 32434 9000 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 11200 0 11400 200 4 DVSS:
port 49 nsew
rlabel metal3 s 11200 32434 11400 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 13600 0 13800 200 4 DVSS:
port 49 nsew
rlabel metal3 s 13600 32434 13800 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 16000 0 16200 200 4 DVSS:
port 49 nsew
rlabel metal3 s 16000 32434 16200 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 18400 0 18600 200 4 DVSS:
port 49 nsew
rlabel metal3 s 18400 32434 18600 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 20800 0 21000 200 4 DVSS:
port 49 nsew
rlabel metal3 s 20800 32434 21000 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 23200 0 23400 200 4 DVSS:
port 49 nsew
rlabel metal3 s 23200 32434 23400 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 25600 0 25800 200 4 DVSS:
port 49 nsew
rlabel metal3 s 25600 32434 25800 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 28000 0 28200 200 4 DVSS:
port 49 nsew
rlabel metal3 s 28000 32434 28200 32634 4 DVSS:
port 49 nsew
rlabel metal3 s 30400 0 30600 200 4 DVSS:
port 49 nsew
rlabel metal3 s 30400 32434 30600 32634 4 DVSS:
port 49 nsew
rlabel metal1 s 0 -49 98 49 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 -49 32064 49 4 DVSS:
port 49 nsew
rlabel metal1 s 0 1283 98 1381 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 1283 32064 1381 4 DVSS:
port 49 nsew
rlabel metal1 s 0 2615 98 2713 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 2615 32064 2713 4 DVSS:
port 49 nsew
rlabel metal1 s 0 3947 98 4045 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 3947 32064 4045 4 DVSS:
port 49 nsew
rlabel metal1 s 0 5279 98 5377 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 5279 32064 5377 4 DVSS:
port 49 nsew
rlabel metal1 s 0 6611 98 6709 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 6611 32064 6709 4 DVSS:
port 49 nsew
rlabel metal1 s 0 7943 98 8041 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 7943 32064 8041 4 DVSS:
port 49 nsew
rlabel metal1 s 0 9275 98 9373 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 9275 32064 9373 4 DVSS:
port 49 nsew
rlabel metal1 s 0 10607 98 10705 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 10607 32064 10705 4 DVSS:
port 49 nsew
rlabel metal1 s 0 11939 98 12037 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 11939 32064 12037 4 DVSS:
port 49 nsew
rlabel metal1 s 0 13271 98 13369 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 13271 32064 13369 4 DVSS:
port 49 nsew
rlabel metal1 s 0 14603 98 14701 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 14603 32064 14701 4 DVSS:
port 49 nsew
rlabel metal1 s 0 15935 98 16033 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 15935 32064 16033 4 DVSS:
port 49 nsew
rlabel metal1 s 0 17267 98 17365 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 17267 32064 17365 4 DVSS:
port 49 nsew
rlabel metal1 s 0 18599 98 18697 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 18599 32064 18697 4 DVSS:
port 49 nsew
rlabel metal1 s 0 19931 98 20029 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 19931 32064 20029 4 DVSS:
port 49 nsew
rlabel metal1 s 0 21263 98 21361 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 21263 32064 21361 4 DVSS:
port 49 nsew
rlabel metal1 s 0 22595 98 22693 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 22595 32064 22693 4 DVSS:
port 49 nsew
rlabel metal1 s 0 23927 98 24025 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 23927 32064 24025 4 DVSS:
port 49 nsew
rlabel metal1 s 0 25259 98 25357 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 25259 32064 25357 4 DVSS:
port 49 nsew
rlabel metal1 s 0 26591 98 26689 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 26591 32064 26689 4 DVSS:
port 49 nsew
rlabel metal1 s 0 27923 98 28021 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 27923 32064 28021 4 DVSS:
port 49 nsew
rlabel metal1 s 0 29255 98 29353 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 29255 32064 29353 4 DVSS:
port 49 nsew
rlabel metal1 s 0 30587 98 30685 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 30587 32064 30685 4 DVSS:
port 49 nsew
rlabel metal1 s 0 31919 98 32017 4 DVSS:
port 49 nsew
rlabel metal1 s 31966 31919 32064 32017 4 DVSS:
port 49 nsew
rlabel metal3 s 400 0 600 200 4 DVDD:
port 50 nsew
rlabel metal3 s 400 32434 600 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 2800 0 3000 200 4 DVDD:
port 50 nsew
rlabel metal3 s 2800 32434 3000 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 5200 0 5400 200 4 DVDD:
port 50 nsew
rlabel metal3 s 5200 32434 5400 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 7600 0 7800 200 4 DVDD:
port 50 nsew
rlabel metal3 s 7600 32434 7800 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 10000 0 10200 200 4 DVDD:
port 50 nsew
rlabel metal3 s 10000 32434 10200 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 12400 0 12600 200 4 DVDD:
port 50 nsew
rlabel metal3 s 12400 32434 12600 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 14800 0 15000 200 4 DVDD:
port 50 nsew
rlabel metal3 s 14800 32434 15000 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 17200 0 17400 200 4 DVDD:
port 50 nsew
rlabel metal3 s 17200 32434 17400 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 19600 0 19800 200 4 DVDD:
port 50 nsew
rlabel metal3 s 19600 32434 19800 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 22000 0 22200 200 4 DVDD:
port 50 nsew
rlabel metal3 s 22000 32434 22200 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 24400 0 24600 200 4 DVDD:
port 50 nsew
rlabel metal3 s 24400 32434 24600 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 26800 0 27000 200 4 DVDD:
port 50 nsew
rlabel metal3 s 26800 32434 27000 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 29200 0 29400 200 4 DVDD:
port 50 nsew
rlabel metal3 s 29200 32434 29400 32634 4 DVDD:
port 50 nsew
rlabel metal3 s 31600 0 31800 200 4 DVDD:
port 50 nsew
rlabel metal3 s 31600 32434 31800 32634 4 DVDD:
port 50 nsew
rlabel metal1 s 0 617 98 715 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 617 32064 715 4 DVDD:
port 50 nsew
rlabel metal1 s 0 1949 98 2047 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 1949 32064 2047 4 DVDD:
port 50 nsew
rlabel metal1 s 0 3281 98 3379 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 3281 32064 3379 4 DVDD:
port 50 nsew
rlabel metal1 s 0 4613 98 4711 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 4613 32064 4711 4 DVDD:
port 50 nsew
rlabel metal1 s 0 5945 98 6043 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 5945 32064 6043 4 DVDD:
port 50 nsew
rlabel metal1 s 0 7277 98 7375 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 7277 32064 7375 4 DVDD:
port 50 nsew
rlabel metal1 s 0 8609 98 8707 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 8609 32064 8707 4 DVDD:
port 50 nsew
rlabel metal1 s 0 9941 98 10039 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 9941 32064 10039 4 DVDD:
port 50 nsew
rlabel metal1 s 0 11273 98 11371 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 11273 32064 11371 4 DVDD:
port 50 nsew
rlabel metal1 s 0 12605 98 12703 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 12605 32064 12703 4 DVDD:
port 50 nsew
rlabel metal1 s 0 13937 98 14035 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 13937 32064 14035 4 DVDD:
port 50 nsew
rlabel metal1 s 0 15269 98 15367 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 15269 32064 15367 4 DVDD:
port 50 nsew
rlabel metal1 s 0 16601 98 16699 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 16601 32064 16699 4 DVDD:
port 50 nsew
rlabel metal1 s 0 17933 98 18031 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 17933 32064 18031 4 DVDD:
port 50 nsew
rlabel metal1 s 0 19265 98 19363 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 19265 32064 19363 4 DVDD:
port 50 nsew
rlabel metal1 s 0 20597 98 20695 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 20597 32064 20695 4 DVDD:
port 50 nsew
rlabel metal1 s 0 21929 98 22027 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 21929 32064 22027 4 DVDD:
port 50 nsew
rlabel metal1 s 0 23261 98 23359 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 23261 32064 23359 4 DVDD:
port 50 nsew
rlabel metal1 s 0 24593 98 24691 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 24593 32064 24691 4 DVDD:
port 50 nsew
rlabel metal1 s 0 25925 98 26023 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 25925 32064 26023 4 DVDD:
port 50 nsew
rlabel metal1 s 0 27257 98 27355 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 27257 32064 27355 4 DVDD:
port 50 nsew
rlabel metal1 s 0 28589 98 28687 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 28589 32064 28687 4 DVDD:
port 50 nsew
rlabel metal1 s 0 29921 98 30019 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 29921 32064 30019 4 DVDD:
port 50 nsew
rlabel metal1 s 0 31253 98 31351 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 31253 32064 31351 4 DVDD:
port 50 nsew
rlabel metal1 s 0 32585 98 32683 4 DVDD:
port 50 nsew
rlabel metal1 s 31966 32585 32064 32683 4 DVDD:
port 50 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 51 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 52 nsew
rlabel metal2 s 48 17649 48 17649 4 clk_out
port 1 nsew
rlabel metal2 s 48 37 48 37 4 div_ratio_half[5]
port 2 nsew
rlabel metal2 s 48 1369 48 1369 4 div_ratio_half[4]
port 3 nsew
rlabel metal2 s 48 2701 48 2701 4 div_ratio_half[3]
port 4 nsew
rlabel metal2 s 48 4107 48 4107 4 div_ratio_half[2]
port 5 nsew
rlabel metal2 s 48 5439 48 5439 4 div_ratio_half[1]
port 6 nsew
rlabel metal2 s 48 6771 48 6771 4 div_ratio_half[0]
port 7 nsew
rlabel metal2 s 48 16317 48 16317 4 ref_clk
port 8 nsew
rlabel metal2 s 48 8103 48 8103 4 rst
port 9 nsew
rlabel metal2 s 48 9509 48 9509 4 aux_osc_en
port 10 nsew
rlabel metal2 s 48 10841 48 10841 4 fftl_en
port 11 nsew
rlabel metal2 s 48 12247 48 12247 4 fine_control_avg_window_select[4]
port 12 nsew
rlabel metal2 s 48 13579 48 13579 4 fine_control_avg_window_select[3]
port 13 nsew
rlabel metal2 s 48 18981 48 18981 4 fine_control_avg_window_select[2]
port 14 nsew
rlabel metal2 s 48 20387 48 20387 4 fine_control_avg_window_select[1]
port 15 nsew
rlabel metal2 s 48 21719 48 21719 4 fine_control_avg_window_select[0]
port 16 nsew
rlabel metal2 s 48 23051 48 23051 4 fine_con_step_size[3]
port 17 nsew
rlabel metal2 s 48 24383 48 24383 4 fine_con_step_size[2]
port 18 nsew
rlabel metal2 s 48 25789 48 25789 4 fine_con_step_size[1]
port 19 nsew
rlabel metal2 s 48 27121 48 27121 4 fine_con_step_size[0]
port 20 nsew
rlabel metal2 s 48 28453 48 28453 4 manual_control_osc[12]
port 21 nsew
rlabel metal2 s 48 29859 48 29859 4 manual_control_osc[11]
port 22 nsew
rlabel metal2 s 48 31191 48 31191 4 manual_control_osc[10]
port 23 nsew
rlabel metal2 s 48 32523 48 32523 4 manual_control_osc[9]
port 24 nsew
rlabel metal2 s 32015 32597 32015 32597 4 manual_control_osc[8]
port 25 nsew
rlabel metal2 s 32015 31117 32015 31117 4 manual_control_osc[7]
port 26 nsew
rlabel metal2 s 32015 29637 32015 29637 4 manual_control_osc[6]
port 27 nsew
rlabel metal2 s 32015 28157 32015 28157 4 manual_control_osc[5]
port 28 nsew
rlabel metal2 s 32015 26677 32015 26677 4 manual_control_osc[4]
port 29 nsew
rlabel metal2 s 32015 25197 32015 25197 4 manual_control_osc[3]
port 30 nsew
rlabel metal2 s 32015 23717 32015 23717 4 manual_control_osc[2]
port 31 nsew
rlabel metal2 s 32015 22237 32015 22237 4 manual_control_osc[1]
port 32 nsew
rlabel metal2 s 32015 20757 32015 20757 4 manual_control_osc[0]
port 33 nsew
rlabel metal2 s 48 14911 48 14911 4 aux_clk_out
port 34 nsew
rlabel metal2 s 32015 19277 32015 19277 4 out_star
port 35 nsew
rlabel metal2 s 32015 17797 32015 17797 4 osc_fine_con_final[12]
port 36 nsew
rlabel metal2 s 32015 16317 32015 16317 4 osc_fine_con_final[11]
port 37 nsew
rlabel metal2 s 32015 14837 32015 14837 4 osc_fine_con_final[10]
port 38 nsew
rlabel metal2 s 32015 13357 32015 13357 4 osc_fine_con_final[9]
port 39 nsew
rlabel metal2 s 32015 11877 32015 11877 4 osc_fine_con_final[8]
port 40 nsew
rlabel metal2 s 32015 10397 32015 10397 4 osc_fine_con_final[7]
port 41 nsew
rlabel metal2 s 32015 8917 32015 8917 4 osc_fine_con_final[6]
port 42 nsew
rlabel metal2 s 32015 7437 32015 7437 4 osc_fine_con_final[5]
port 43 nsew
rlabel metal2 s 32015 5957 32015 5957 4 osc_fine_con_final[4]
port 44 nsew
rlabel metal2 s 32015 4477 32015 4477 4 osc_fine_con_final[3]
port 45 nsew
rlabel metal2 s 32015 2997 32015 2997 4 osc_fine_con_final[2]
port 46 nsew
rlabel metal2 s 32015 1517 32015 1517 4 osc_fine_con_final[1]
port 47 nsew
rlabel metal2 s 32015 37 32015 37 4 osc_fine_con_final[0]
port 48 nsew
rlabel metal3 s 1700 100 1700 100 4 DVSS:
port 49 nsew
rlabel metal3 s 1700 32534 1700 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 4100 100 4100 100 4 DVSS:
port 49 nsew
rlabel metal3 s 4100 32534 4100 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 6500 100 6500 100 4 DVSS:
port 49 nsew
rlabel metal3 s 6500 32534 6500 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 8900 100 8900 100 4 DVSS:
port 49 nsew
rlabel metal3 s 8900 32534 8900 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 11300 100 11300 100 4 DVSS:
port 49 nsew
rlabel metal3 s 11300 32534 11300 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 13700 100 13700 100 4 DVSS:
port 49 nsew
rlabel metal3 s 13700 32534 13700 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 16100 100 16100 100 4 DVSS:
port 49 nsew
rlabel metal3 s 16100 32534 16100 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 18500 100 18500 100 4 DVSS:
port 49 nsew
rlabel metal3 s 18500 32534 18500 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 20900 100 20900 100 4 DVSS:
port 49 nsew
rlabel metal3 s 20900 32534 20900 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 23300 100 23300 100 4 DVSS:
port 49 nsew
rlabel metal3 s 23300 32534 23300 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 25700 100 25700 100 4 DVSS:
port 49 nsew
rlabel metal3 s 25700 32534 25700 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 28100 100 28100 100 4 DVSS:
port 49 nsew
rlabel metal3 s 28100 32534 28100 32534 4 DVSS:
port 49 nsew
rlabel metal3 s 30500 100 30500 100 4 DVSS:
port 49 nsew
rlabel metal3 s 30500 32534 30500 32534 4 DVSS:
port 49 nsew
rlabel metal1 s 49 0 49 0 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 0 32015 0 4 DVSS:
port 49 nsew
rlabel metal1 s 49 1332 49 1332 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 1332 32015 1332 4 DVSS:
port 49 nsew
rlabel metal1 s 49 2664 49 2664 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 2664 32015 2664 4 DVSS:
port 49 nsew
rlabel metal1 s 49 3996 49 3996 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 3996 32015 3996 4 DVSS:
port 49 nsew
rlabel metal1 s 49 5328 49 5328 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 5328 32015 5328 4 DVSS:
port 49 nsew
rlabel metal1 s 49 6660 49 6660 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 6660 32015 6660 4 DVSS:
port 49 nsew
rlabel metal1 s 49 7992 49 7992 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 7992 32015 7992 4 DVSS:
port 49 nsew
rlabel metal1 s 49 9324 49 9324 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 9324 32015 9324 4 DVSS:
port 49 nsew
rlabel metal1 s 49 10656 49 10656 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 10656 32015 10656 4 DVSS:
port 49 nsew
rlabel metal1 s 49 11988 49 11988 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 11988 32015 11988 4 DVSS:
port 49 nsew
rlabel metal1 s 49 13320 49 13320 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 13320 32015 13320 4 DVSS:
port 49 nsew
rlabel metal1 s 49 14652 49 14652 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 14652 32015 14652 4 DVSS:
port 49 nsew
rlabel metal1 s 49 15984 49 15984 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 15984 32015 15984 4 DVSS:
port 49 nsew
rlabel metal1 s 49 17316 49 17316 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 17316 32015 17316 4 DVSS:
port 49 nsew
rlabel metal1 s 49 18648 49 18648 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 18648 32015 18648 4 DVSS:
port 49 nsew
rlabel metal1 s 49 19980 49 19980 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 19980 32015 19980 4 DVSS:
port 49 nsew
rlabel metal1 s 49 21312 49 21312 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 21312 32015 21312 4 DVSS:
port 49 nsew
rlabel metal1 s 49 22644 49 22644 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 22644 32015 22644 4 DVSS:
port 49 nsew
rlabel metal1 s 49 23976 49 23976 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 23976 32015 23976 4 DVSS:
port 49 nsew
rlabel metal1 s 49 25308 49 25308 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 25308 32015 25308 4 DVSS:
port 49 nsew
rlabel metal1 s 49 26640 49 26640 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 26640 32015 26640 4 DVSS:
port 49 nsew
rlabel metal1 s 49 27972 49 27972 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 27972 32015 27972 4 DVSS:
port 49 nsew
rlabel metal1 s 49 29304 49 29304 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 29304 32015 29304 4 DVSS:
port 49 nsew
rlabel metal1 s 49 30636 49 30636 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 30636 32015 30636 4 DVSS:
port 49 nsew
rlabel metal1 s 49 31968 49 31968 4 DVSS:
port 49 nsew
rlabel metal1 s 32015 31968 32015 31968 4 DVSS:
port 49 nsew
rlabel metal3 s 500 100 500 100 4 DVDD:
port 50 nsew
rlabel metal3 s 500 32534 500 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 2900 100 2900 100 4 DVDD:
port 50 nsew
rlabel metal3 s 2900 32534 2900 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 5300 100 5300 100 4 DVDD:
port 50 nsew
rlabel metal3 s 5300 32534 5300 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 7700 100 7700 100 4 DVDD:
port 50 nsew
rlabel metal3 s 7700 32534 7700 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 10100 100 10100 100 4 DVDD:
port 50 nsew
rlabel metal3 s 10100 32534 10100 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 12500 100 12500 100 4 DVDD:
port 50 nsew
rlabel metal3 s 12500 32534 12500 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 14900 100 14900 100 4 DVDD:
port 50 nsew
rlabel metal3 s 14900 32534 14900 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 17300 100 17300 100 4 DVDD:
port 50 nsew
rlabel metal3 s 17300 32534 17300 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 19700 100 19700 100 4 DVDD:
port 50 nsew
rlabel metal3 s 19700 32534 19700 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 22100 100 22100 100 4 DVDD:
port 50 nsew
rlabel metal3 s 22100 32534 22100 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 24500 100 24500 100 4 DVDD:
port 50 nsew
rlabel metal3 s 24500 32534 24500 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 26900 100 26900 100 4 DVDD:
port 50 nsew
rlabel metal3 s 26900 32534 26900 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 29300 100 29300 100 4 DVDD:
port 50 nsew
rlabel metal3 s 29300 32534 29300 32534 4 DVDD:
port 50 nsew
rlabel metal3 s 31700 100 31700 100 4 DVDD:
port 50 nsew
rlabel metal3 s 31700 32534 31700 32534 4 DVDD:
port 50 nsew
rlabel metal1 s 49 666 49 666 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 666 32015 666 4 DVDD:
port 50 nsew
rlabel metal1 s 49 1998 49 1998 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 1998 32015 1998 4 DVDD:
port 50 nsew
rlabel metal1 s 49 3330 49 3330 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 3330 32015 3330 4 DVDD:
port 50 nsew
rlabel metal1 s 49 4662 49 4662 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 4662 32015 4662 4 DVDD:
port 50 nsew
rlabel metal1 s 49 5994 49 5994 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 5994 32015 5994 4 DVDD:
port 50 nsew
rlabel metal1 s 49 7326 49 7326 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 7326 32015 7326 4 DVDD:
port 50 nsew
rlabel metal1 s 49 8658 49 8658 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 8658 32015 8658 4 DVDD:
port 50 nsew
rlabel metal1 s 49 9990 49 9990 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 9990 32015 9990 4 DVDD:
port 50 nsew
rlabel metal1 s 49 11322 49 11322 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 11322 32015 11322 4 DVDD:
port 50 nsew
rlabel metal1 s 49 12654 49 12654 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 12654 32015 12654 4 DVDD:
port 50 nsew
rlabel metal1 s 49 13986 49 13986 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 13986 32015 13986 4 DVDD:
port 50 nsew
rlabel metal1 s 49 15318 49 15318 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 15318 32015 15318 4 DVDD:
port 50 nsew
rlabel metal1 s 49 16650 49 16650 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 16650 32015 16650 4 DVDD:
port 50 nsew
rlabel metal1 s 49 17982 49 17982 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 17982 32015 17982 4 DVDD:
port 50 nsew
rlabel metal1 s 49 19314 49 19314 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 19314 32015 19314 4 DVDD:
port 50 nsew
rlabel metal1 s 49 20646 49 20646 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 20646 32015 20646 4 DVDD:
port 50 nsew
rlabel metal1 s 49 21978 49 21978 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 21978 32015 21978 4 DVDD:
port 50 nsew
rlabel metal1 s 49 23310 49 23310 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 23310 32015 23310 4 DVDD:
port 50 nsew
rlabel metal1 s 49 24642 49 24642 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 24642 32015 24642 4 DVDD:
port 50 nsew
rlabel metal1 s 49 25974 49 25974 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 25974 32015 25974 4 DVDD:
port 50 nsew
rlabel metal1 s 49 27306 49 27306 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 27306 32015 27306 4 DVDD:
port 50 nsew
rlabel metal1 s 49 28638 49 28638 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 28638 32015 28638 4 DVDD:
port 50 nsew
rlabel metal1 s 49 29970 49 29970 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 29970 32015 29970 4 DVDD:
port 50 nsew
rlabel metal1 s 49 31302 49 31302 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 31302 32015 31302 4 DVDD:
port 50 nsew
rlabel metal1 s 49 32634 49 32634 4 DVDD:
port 50 nsew
rlabel metal1 s 32015 32634 32015 32634 4 DVDD:
port 50 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 51 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 52 nsew
<< properties >>
string path 498.000 541.125 502.800 541.125 
<< end >>
