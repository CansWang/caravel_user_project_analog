magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal2 >>
rect -139 28 139 33
rect -139 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 139 28
rect -139 -33 139 -28
<< via2 >>
rect -108 -28 -52 28
rect -28 -28 28 28
rect 52 -28 108 28
<< metal3 >>
rect -139 28 139 33
rect -139 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 139 28
rect -139 -33 139 -28
<< end >>
