magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal2 >>
rect -100 28 100 49
rect -100 -28 -68 28
rect -12 -28 12 28
rect 68 -28 100 28
rect -100 -49 100 -28
<< via2 >>
rect -68 -28 -12 28
rect 12 -28 68 28
<< metal3 >>
rect -100 28 100 49
rect -100 -28 -68 28
rect -12 -28 12 28
rect 68 -28 100 28
rect -100 -49 100 -28
<< end >>
