magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< error_s >>
rect 1118 9435 1119 9480
rect 2366 9435 2367 9480
rect 3710 9435 3711 9480
rect 4574 9435 4575 9480
rect 5534 9435 5535 9480
rect 6782 9435 6783 9480
rect 8030 9435 8031 9480
rect 9278 9435 9279 9480
rect 350 9179 351 9224
rect 1790 9179 1791 9224
rect 5534 9179 5535 9224
rect 6782 9179 6783 9224
rect 8030 9179 8031 9224
rect 9374 9179 9375 9224
rect 5534 8103 5535 8148
rect 6782 8103 6783 8148
rect 8030 8103 8031 8148
rect 9278 8103 9279 8148
rect 1790 7847 1791 7892
rect 6782 7847 6783 7892
rect 8030 7847 8031 7892
rect 9374 7847 9375 7892
rect 5534 6771 5535 6816
rect 8702 6771 8703 6816
rect 4094 6515 4095 6560
rect 8030 6515 8031 6560
rect 9374 6515 9375 6560
rect 4574 5439 4575 5484
rect 5534 5183 5535 5228
rect 6782 5183 6783 5228
rect 8030 5183 8031 5228
rect 2366 4107 2367 4152
rect 5534 4107 5535 4152
rect 9566 3851 9567 3896
rect 9278 2775 9279 2820
rect 9374 2519 9375 2564
rect 6206 1443 6207 1488
rect 7262 1443 7263 1488
rect 9374 1187 9375 1232
rect 6206 111 6207 156
rect 7070 111 7071 156
rect 8030 111 8031 156
rect 9278 111 9279 156
<< locali >>
rect 3871 8120 3905 8564
rect 3967 8342 4001 8564
rect 3967 8308 4080 8342
rect 3871 8086 4080 8120
rect 4543 7642 4656 7676
rect 4543 7420 4577 7642
rect 5232 7420 5345 7454
rect 3775 4346 3809 4494
rect 3696 4312 3809 4346
rect 6079 3498 6113 3902
rect 4560 982 4848 1016
<< metal1 >>
rect 0 10607 10080 10705
rect 322 10235 3614 10263
rect 322 10115 350 10235
rect 130 10087 350 10115
rect 3586 10115 3614 10235
rect 3586 10087 3806 10115
rect 0 9941 10080 10039
rect 34 9717 3230 9745
rect 3033 9421 3120 9449
rect 0 9275 10080 9373
rect 130 9051 1022 9079
rect 3010 9051 3134 9079
rect 2553 8977 2640 9005
rect 4546 8977 4670 9005
rect 802 8903 926 8931
rect 4089 8755 4176 8783
rect 4665 8755 4752 8783
rect 0 8609 10080 8707
rect 34 8533 446 8561
rect 2146 8533 3902 8561
rect 3970 8533 4190 8561
rect 418 8487 446 8533
rect 418 8459 926 8487
rect 2914 8459 4478 8487
rect 898 8413 926 8459
rect 898 8385 2078 8413
rect 2050 8339 2078 8385
rect 2722 8385 3422 8413
rect 2722 8339 2750 8385
rect 322 8311 446 8339
rect 729 8311 816 8339
rect 2050 8311 2750 8339
rect 2928 8311 3015 8339
rect 3106 8311 4190 8339
rect 4326 8191 4354 8339
rect 4450 8321 4478 8459
rect 4326 8163 4766 8191
rect 3225 8089 3312 8117
rect 4642 8089 4958 8117
rect 0 7943 10080 8041
rect 4354 7867 4670 7895
rect 34 7747 62 7821
rect 4834 7793 5726 7821
rect 34 7719 1118 7747
rect 3010 7719 3326 7747
rect 5026 7691 5054 7747
rect 2553 7645 2640 7673
rect 4812 7645 4916 7673
rect 5122 7645 5630 7673
rect 5122 7599 5150 7645
rect 537 7571 624 7599
rect 706 7525 734 7599
rect 898 7571 1022 7599
rect 3490 7571 4382 7599
rect 4546 7571 5150 7599
rect 3490 7525 3518 7571
rect 130 7497 734 7525
rect 2338 7497 3518 7525
rect 2338 7451 2366 7497
rect 2146 7423 2366 7451
rect 4354 7451 4382 7571
rect 5794 7497 6302 7525
rect 5794 7451 5822 7497
rect 4354 7423 4574 7451
rect 5314 7423 5822 7451
rect 6274 7451 6302 7497
rect 6274 7423 6494 7451
rect 0 7277 10080 7375
rect 2073 7201 2160 7229
rect 34 7127 1118 7155
rect 1090 7081 1118 7127
rect 2146 7127 2942 7155
rect 2146 7081 2174 7127
rect 1090 7053 2174 7081
rect 4642 7053 4766 7081
rect 322 6979 446 7007
rect 802 6979 926 7007
rect 2338 6979 2654 7007
rect 4546 6979 4862 7007
rect 5602 6979 6398 7007
rect 6466 6979 6782 7007
rect 2722 6905 3326 6933
rect 3298 6831 3326 6905
rect 4066 6757 4286 6785
rect 7522 6757 7934 6785
rect 0 6611 10080 6709
rect 2818 6535 3134 6563
rect 3202 6535 3326 6563
rect 514 6387 734 6415
rect 2841 6387 2928 6415
rect 4930 6387 6014 6415
rect 130 6313 350 6341
rect 4546 6313 4670 6341
rect 5529 6313 5616 6341
rect 226 6239 3326 6267
rect 1785 6091 1872 6119
rect 4834 6091 5150 6119
rect 7257 6091 7344 6119
rect 0 5945 10080 6043
rect 4066 5721 4670 5749
rect 4642 5675 4670 5721
rect 322 5647 446 5675
rect 2338 5647 2654 5675
rect 2722 5647 3134 5675
rect 4642 5647 5150 5675
rect 5218 5647 5438 5675
rect 5506 5601 5534 5675
rect 5602 5647 5822 5675
rect 7714 5647 7934 5675
rect 802 5573 1022 5601
rect 5314 5573 5534 5601
rect 6105 5573 6192 5601
rect 6370 5573 8126 5601
rect 6370 5527 6398 5573
rect 4450 5499 4958 5527
rect 5698 5499 6398 5527
rect 8578 5499 9086 5527
rect 4450 5453 4478 5499
rect 2073 5425 2160 5453
rect 4258 5425 4478 5453
rect 4930 5453 4958 5499
rect 8578 5453 8606 5499
rect 4930 5425 5150 5453
rect 7522 5425 8126 5453
rect 8386 5425 8606 5453
rect 9058 5453 9086 5499
rect 9058 5425 9278 5453
rect 0 5279 10080 5377
rect 1858 5203 2654 5231
rect 3202 5203 3422 5231
rect 3394 5194 3422 5203
rect 5986 5203 6206 5231
rect 3394 5166 5534 5194
rect 5506 5157 5534 5166
rect 5986 5157 6014 5203
rect 5506 5129 6014 5157
rect 4450 5055 5342 5083
rect 130 4981 350 5009
rect 514 4981 734 5009
rect 2146 4981 2654 5009
rect 2914 4935 2942 5009
rect 3010 4981 3326 5009
rect 3874 4981 4670 5009
rect 4834 4935 4862 5009
rect 8290 4981 9086 5009
rect 8290 4935 8318 4981
rect 2914 4907 3710 4935
rect 3778 4907 3998 4935
rect 3970 4861 3998 4907
rect 4642 4907 8318 4935
rect 4642 4861 4670 4907
rect 3970 4833 4670 4861
rect 898 4759 1694 4787
rect 4953 4759 5040 4787
rect 8770 4759 9086 4787
rect 0 4613 10080 4711
rect 3778 4463 4574 4491
rect 9442 4463 10046 4491
rect 322 4389 2654 4417
rect 3298 4389 3518 4417
rect 34 4315 734 4343
rect 3874 4315 4286 4343
rect 8866 4315 9854 4343
rect 226 4241 1118 4269
rect 1762 4241 3038 4269
rect 9154 4241 9278 4269
rect 610 4093 734 4121
rect 921 4093 1008 4121
rect 4450 4093 4766 4121
rect 6946 4093 7742 4121
rect 0 3947 10080 4045
rect 34 3871 542 3899
rect 6082 3871 6782 3899
rect 7330 3871 7454 3899
rect 7906 3871 8798 3899
rect 514 3825 542 3871
rect 7906 3825 7934 3871
rect 514 3797 1406 3825
rect 6178 3797 7934 3825
rect 1378 3751 1406 3797
rect 1378 3723 2270 3751
rect 4738 3723 5822 3751
rect 130 3649 350 3677
rect 514 3649 734 3677
rect 706 3603 734 3649
rect 1186 3649 1598 3677
rect 3129 3649 3216 3677
rect 5410 3649 6302 3677
rect 1186 3603 1214 3649
rect 706 3575 1214 3603
rect 1570 3603 1598 3649
rect 6352 3640 6416 3763
rect 8770 3751 8798 3871
rect 9538 3871 9758 3899
rect 9538 3751 9566 3871
rect 7522 3677 7550 3751
rect 7714 3723 8222 3751
rect 8770 3723 9566 3751
rect 6466 3603 6494 3677
rect 6681 3649 6768 3677
rect 6969 3649 7056 3677
rect 7138 3649 7262 3677
rect 7426 3649 7550 3677
rect 8194 3677 8222 3723
rect 8194 3649 8606 3677
rect 7138 3603 7166 3649
rect 1570 3575 2174 3603
rect 6466 3575 7166 3603
rect 7833 3575 7920 3603
rect 6082 3501 6686 3529
rect 6850 3501 7070 3529
rect 1378 3427 1694 3455
rect 6274 3427 8702 3455
rect 0 3281 10080 3379
rect 8098 3205 8606 3233
rect 8578 3159 8606 3205
rect 9826 3205 10046 3233
rect 9826 3159 9854 3205
rect 8578 3131 9854 3159
rect 1090 3057 3600 3085
rect 7426 3057 8414 3085
rect 1090 3011 1118 3057
rect 7426 3011 7454 3057
rect 130 2983 1118 3011
rect 1200 2983 1287 3011
rect 3129 2983 3216 3011
rect 5529 2983 5616 3011
rect 7234 2983 7454 3011
rect 610 2909 926 2937
rect 1570 2909 2174 2937
rect 4834 2909 6014 2937
rect 4834 2863 4862 2909
rect 3394 2835 3998 2863
rect 3970 2826 3998 2835
rect 4642 2835 4862 2863
rect 4642 2826 4670 2835
rect 3970 2798 4670 2826
rect 7234 2789 7262 2983
rect 7522 2937 7550 3011
rect 7618 2983 7838 3011
rect 7920 2983 8007 3011
rect 8217 2983 8304 3011
rect 8409 2983 8496 3011
rect 8592 2983 8679 3011
rect 8770 2983 9470 3011
rect 7522 2909 8126 2937
rect 7330 2835 7646 2863
rect 7618 2789 7646 2835
rect 34 2761 734 2789
rect 2914 2761 3806 2789
rect 7234 2761 7550 2789
rect 7618 2761 8222 2789
rect 0 2615 10080 2713
rect 825 2539 912 2567
rect 2073 2539 2160 2567
rect 6658 2539 7070 2567
rect 7618 2539 8510 2567
rect 1090 2502 1886 2530
rect 1090 2493 1118 2502
rect 226 2465 1118 2493
rect 1858 2493 1886 2502
rect 1858 2465 2270 2493
rect 802 2391 1982 2419
rect 2242 2391 2270 2465
rect 3010 2391 3134 2419
rect 802 2345 830 2391
rect 441 2317 528 2345
rect 610 2317 830 2345
rect 898 2317 1406 2345
rect 1858 2317 2462 2345
rect 2553 2317 2640 2345
rect 3202 2317 4574 2345
rect 5506 2317 5630 2345
rect 5794 2317 5918 2345
rect 8482 2317 8702 2345
rect 2434 2271 2462 2317
rect 3202 2271 3230 2317
rect 34 2243 638 2271
rect 1017 2243 1104 2271
rect 610 2197 638 2243
rect 1186 2197 1214 2271
rect 2434 2243 3230 2271
rect 4665 2243 4752 2271
rect 610 2169 1214 2197
rect 1378 2132 2270 2160
rect 1378 2123 1406 2132
rect 322 2095 1406 2123
rect 2242 2123 2270 2132
rect 2242 2095 3422 2123
rect 4354 2095 5150 2123
rect 0 1949 10080 2047
rect 3010 1873 3518 1901
rect 3490 1864 3518 1873
rect 5602 1873 5822 1901
rect 8290 1873 8510 1901
rect 5602 1864 5630 1873
rect 3490 1836 5630 1864
rect 8482 1827 8510 1873
rect 9058 1873 9278 1901
rect 9058 1827 9086 1873
rect 706 1799 3326 1827
rect 8482 1799 9086 1827
rect 3106 1725 3230 1753
rect 3298 1725 3326 1799
rect 4642 1725 5246 1753
rect 5218 1679 5246 1725
rect 322 1651 446 1679
rect 802 1651 1118 1679
rect 1858 1651 2462 1679
rect 2722 1531 2750 1679
rect 2818 1651 2942 1679
rect 3874 1651 4574 1679
rect 5049 1651 5136 1679
rect 5218 1651 5438 1679
rect 5506 1605 5534 1679
rect 7714 1651 7934 1679
rect 4738 1577 5534 1605
rect 5698 1577 8126 1605
rect 2722 1503 3710 1531
rect 3970 1466 4958 1494
rect 3970 1457 3998 1466
rect 2146 1429 2462 1457
rect 3778 1429 3998 1457
rect 4930 1457 4958 1466
rect 4930 1429 5150 1457
rect 0 1283 10080 1381
rect 34 1207 542 1235
rect 1785 1207 1872 1235
rect 6850 1207 7166 1235
rect 8482 1207 9182 1235
rect 514 1161 542 1207
rect 514 1133 1694 1161
rect 1666 1087 1694 1133
rect 1666 1059 2270 1087
rect 2914 1059 3806 1087
rect 130 985 350 1013
rect 514 985 1598 1013
rect 3970 985 4574 1013
rect 5529 985 5616 1013
rect 5794 985 6014 1013
rect 7906 985 8222 1013
rect 1570 939 1598 985
rect 1570 911 2174 939
rect 2434 911 2750 939
rect 514 837 1406 865
rect 514 791 542 837
rect 1378 828 1406 837
rect 1378 800 2654 828
rect 34 763 542 791
rect 2626 791 2654 800
rect 2818 791 2846 939
rect 3033 911 3120 939
rect 3202 911 3326 939
rect 4354 911 5534 939
rect 2626 763 2846 791
rect 5049 763 5136 791
rect 0 617 10080 715
rect 5698 541 5822 569
rect 34 467 3326 495
rect 4354 393 4766 421
rect 4738 347 4766 393
rect 322 319 446 347
rect 802 319 1022 347
rect 994 273 1022 319
rect 1954 319 2462 347
rect 2553 319 2640 347
rect 3010 319 3134 347
rect 4738 319 5150 347
rect 5218 319 5438 347
rect 5520 319 5607 347
rect 1954 273 1982 319
rect 994 245 1982 273
rect 3298 245 4190 273
rect 3298 199 3326 245
rect 2338 171 3326 199
rect 4162 199 4190 245
rect 7234 245 9854 273
rect 7234 199 7262 245
rect 4162 171 4574 199
rect 7042 171 7262 199
rect 9826 199 9854 245
rect 9826 171 10046 199
rect 2338 125 2366 171
rect 2146 97 2366 125
rect 4546 125 4574 171
rect 4546 97 5150 125
rect 0 -49 10080 49
<< metal2 >>
rect 0 10605 97 10633
rect 34 9967 62 10605
rect 130 10087 158 10656
rect 9730 10605 10080 10633
rect 34 9939 158 9967
rect 0 9865 97 9893
rect 34 9717 62 9865
rect 0 9125 97 9153
rect 34 8533 62 9125
rect 130 9051 158 9939
rect 3106 9051 3134 9449
rect 0 8459 97 8487
rect 34 7793 62 8459
rect 0 7719 97 7747
rect 34 7599 62 7719
rect 34 7571 254 7599
rect 34 7081 62 7155
rect 0 7053 97 7081
rect 130 6341 158 7525
rect 0 6313 158 6341
rect 226 6239 254 7571
rect 0 5647 97 5675
rect 34 5009 62 5647
rect 34 4981 158 5009
rect 0 4907 97 4935
rect 34 4315 62 4907
rect 130 4343 158 4981
rect 130 4315 254 4343
rect 0 4241 97 4269
rect 226 4241 254 4315
rect 34 3871 62 4241
rect 0 3501 97 3529
rect 34 3085 62 3501
rect 34 3057 254 3085
rect 0 2835 97 2863
rect 34 2761 62 2835
rect 34 2123 62 2271
rect 0 2095 97 2123
rect 0 1429 97 1457
rect 34 1207 62 1429
rect 34 717 62 791
rect 0 689 97 717
rect 34 51 62 495
rect 0 23 97 51
rect 130 0 158 3011
rect 226 2465 254 3057
rect 322 319 350 8339
rect 802 8311 830 8931
rect 610 7451 638 7599
rect 610 7423 734 7451
rect 706 6387 734 7423
rect 898 6979 926 7599
rect 2146 7201 2174 7451
rect 706 4093 734 5009
rect 898 4639 926 4787
rect 850 4611 926 4639
rect 850 4047 878 4611
rect 994 4093 1022 5601
rect 1858 5203 1886 6119
rect 2146 4981 2174 5453
rect 850 4019 926 4047
rect 610 2715 638 2937
rect 514 2687 638 2715
rect 514 2317 542 2687
rect 706 1799 734 2789
rect 898 2539 926 4019
rect 1186 2983 1214 4417
rect 1378 2317 1406 3455
rect 2146 2539 2174 2937
rect 1090 1651 1118 2271
rect 1858 1207 1886 1679
rect 2434 319 2462 939
rect 2626 319 2654 9005
rect 2914 8311 2942 8487
rect 3298 7719 3326 8117
rect 2914 6387 2942 7155
rect 3106 5647 3134 6563
rect 3298 6535 3326 6859
rect 3298 4389 3326 5009
rect 3778 4907 3806 10115
rect 4162 8533 4190 8783
rect 4546 8339 4574 9005
rect 4162 8311 4574 8339
rect 4258 5425 4286 6785
rect 3010 4047 3038 4269
rect 3202 4047 3230 4199
rect 3874 4171 3902 4343
rect 3010 4019 3230 4047
rect 3202 2983 3230 4019
rect 3106 1725 3134 2419
rect 3394 2095 3422 2863
rect 2914 1059 2942 1679
rect 3778 1429 3806 2789
rect 4546 985 4574 8311
rect 4738 8163 4766 8783
rect 4834 7645 4862 7821
rect 4738 7053 4766 7615
rect 4930 6387 4958 8117
rect 5026 7587 5054 7747
rect 5122 5897 5150 6119
rect 5122 5869 5246 5897
rect 5218 5647 5246 5869
rect 5314 5055 5342 5601
rect 4738 3723 4766 4121
rect 5026 3575 5054 4787
rect 5602 3751 5630 7007
rect 6466 6979 6494 7451
rect 7330 5971 7358 6119
rect 7234 5943 7358 5971
rect 6178 5203 6206 5601
rect 7234 4047 7262 5943
rect 7234 4019 7358 4047
rect 7330 3871 7358 4019
rect 5602 3723 7454 3751
rect 7522 3723 7550 6785
rect 7714 3723 7742 4121
rect 4738 1577 4766 2271
rect 5122 1651 5150 2123
rect 5602 985 5630 3723
rect 6274 3427 6302 3677
rect 6754 3529 6782 3677
rect 7042 3649 7070 3723
rect 7426 3677 7454 3723
rect 7906 3677 7934 5675
rect 6658 2539 6686 3529
rect 6754 3501 6878 3529
rect 6850 2419 6878 3501
rect 6754 2391 6878 2419
rect 5794 1873 5822 2345
rect 6754 1531 6782 2391
rect 6754 1503 6878 1531
rect 6850 1207 6878 1503
rect 3106 319 3134 939
rect 3298 467 3326 939
rect 5122 569 5150 791
rect 5122 541 5246 569
rect 5218 319 5246 541
rect 5506 319 5534 939
rect 5794 541 5822 1013
rect 7042 171 7070 3529
rect 7234 2567 7262 3677
rect 7426 3649 7934 3677
rect 7618 2567 7646 3011
rect 7234 2539 7646 2567
rect 7906 985 7934 3649
rect 8098 2909 8126 5453
rect 8386 3057 8414 5453
rect 8770 4389 8798 4787
rect 8290 1873 8318 3011
rect 8482 2539 8510 3011
rect 8578 2951 8606 3011
rect 8674 2317 8702 3455
rect 9154 1207 9182 4269
rect 9442 2983 9470 4491
rect 9730 3871 9758 10605
rect 9983 7127 10080 7155
rect 10018 4463 10046 7127
rect 9826 4315 9950 4343
rect 9922 0 9950 4315
rect 9983 3575 10080 3603
rect 10018 3205 10046 3575
rect 10018 51 10046 199
rect 9983 23 10080 51
<< metal3 >>
rect 400 0 600 10656
rect 1600 0 1800 10656
rect 2800 0 3000 10656
rect 3186 4155 3918 4215
rect 4000 0 4200 10656
rect 4722 7571 5070 7631
rect 5200 0 5400 10656
rect 6400 0 6600 10656
rect 7600 0 7800 10656
rect 7890 2935 8622 2995
rect 8800 0 9000 10656
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_18
timestamp 1626908933
transform 1 0 0 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_79
timestamp 1626908933
transform 1 0 0 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_64
timestamp 1626908933
transform 1 0 192 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_66
timestamp 1626908933
transform 1 0 0 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_183
timestamp 1626908933
transform 1 0 192 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_185
timestamp 1626908933
transform 1 0 0 0 -1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_179
timestamp 1626908933
transform 1 0 48 0 1 481
box -32 -32 32 32
use M1M2_PR  M1M2_PR_379
timestamp 1626908933
transform 1 0 48 0 1 481
box -32 -32 32 32
use L1M1_PR  L1M1_PR_340
timestamp 1626908933
transform 1 0 432 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_120
timestamp 1626908933
transform 1 0 432 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_300
timestamp 1626908933
transform 1 0 336 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_100
timestamp 1626908933
transform 1 0 336 0 1 333
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_91
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_31
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_91
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_31
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_89
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_44
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use L1M1_PR  L1M1_PR_163
timestamp 1626908933
transform 1 0 816 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_383
timestamp 1626908933
transform 1 0 816 0 1 333
box -29 -23 29 23
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_7
timestamp 1626908933
transform 1 0 1700 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_15
timestamp 1626908933
transform 1 0 1700 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_7
timestamp 1626908933
transform 1 0 1700 0 1 23
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_15
timestamp 1626908933
transform 1 0 1700 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_19
timestamp 1626908933
transform 1 0 2016 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_3
timestamp 1626908933
transform 1 0 2016 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_19
timestamp 1626908933
transform 1 0 2304 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_80
timestamp 1626908933
transform 1 0 2304 0 1 0
box -38 -49 230 715
use L1M1_PR  L1M1_PR_103
timestamp 1626908933
transform 1 0 2160 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_323
timestamp 1626908933
transform 1 0 2160 0 1 111
box -29 -23 29 23
use M1M2_PR  M1M2_PR_335
timestamp 1626908933
transform 1 0 2448 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_135
timestamp 1626908933
transform 1 0 2448 0 1 333
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_186
timestamp 1626908933
transform 1 0 2400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_67
timestamp 1626908933
transform 1 0 2400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_88
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_84
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_43
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_39
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_331
timestamp 1626908933
transform 1 0 2640 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_111
timestamp 1626908933
transform 1 0 2640 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_288
timestamp 1626908933
transform 1 0 2640 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_88
timestamp 1626908933
transform 1 0 2640 0 1 333
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_6
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_22
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_40
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_35
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_28
timestamp 1626908933
transform 1 0 96 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_16
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_11
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_4
timestamp 1626908933
transform 1 0 96 0 -1 1332
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_143
timestamp 1626908933
transform 1 0 3120 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_343
timestamp 1626908933
transform 1 0 3120 0 1 333
box -32 -32 32 32
use L1M1_PR  L1M1_PR_171
timestamp 1626908933
transform 1 0 3024 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_391
timestamp 1626908933
transform 1 0 3024 0 1 333
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_23
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_83
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_23
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_83
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_21
timestamp 1626908933
transform 1 0 3360 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_82
timestamp 1626908933
transform 1 0 3360 0 -1 1332
box -38 -49 230 715
use M1M2_PR  M1M2_PR_178
timestamp 1626908933
transform 1 0 3312 0 1 481
box -32 -32 32 32
use M1M2_PR  M1M2_PR_378
timestamp 1626908933
transform 1 0 3312 0 1 481
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_26
timestamp 1626908933
transform 1 0 2976 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_10
timestamp 1626908933
transform 1 0 2976 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_68
timestamp 1626908933
transform 1 0 4032 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_187
timestamp 1626908933
transform 1 0 4032 0 -1 1332
box -38 -49 134 715
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_6
timestamp 1626908933
transform 1 0 4100 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_14
timestamp 1626908933
transform 1 0 4100 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_6
timestamp 1626908933
transform 1 0 4100 0 1 23
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_14
timestamp 1626908933
transform 1 0 4100 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_15
timestamp 1626908933
transform 1 0 4128 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_13
timestamp 1626908933
transform 1 0 3552 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_7
timestamp 1626908933
transform 1 0 4128 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_5
timestamp 1626908933
transform 1 0 3552 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_22
timestamp 1626908933
transform 1 0 4608 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_83
timestamp 1626908933
transform 1 0 4608 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_63
timestamp 1626908933
transform 1 0 4512 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_182
timestamp 1626908933
transform 1 0 4512 0 1 0
box -38 -49 134 715
use L1M1_PR  L1M1_PR_101
timestamp 1626908933
transform 1 0 4368 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_321
timestamp 1626908933
transform 1 0 4368 0 1 407
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_42
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_87
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_18
timestamp 1626908933
transform 1 0 4800 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_7
timestamp 1626908933
transform 1 0 4800 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_36
timestamp 1626908933
transform 1 0 4608 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_90
timestamp 1626908933
transform 1 0 4608 0 1 0
box -38 -49 422 715
use L1M1_PR  L1M1_PR_322
timestamp 1626908933
transform 1 0 5136 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_320
timestamp 1626908933
transform 1 0 5136 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_102
timestamp 1626908933
transform 1 0 5136 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_100
timestamp 1626908933
transform 1 0 5136 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_242
timestamp 1626908933
transform 1 0 5232 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_42
timestamp 1626908933
transform 1 0 5232 0 1 333
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_75
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_15
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_75
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_15
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_84
timestamp 1626908933
transform 1 0 5280 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_23
timestamp 1626908933
transform 1 0 5280 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_69
timestamp 1626908933
transform 1 0 5472 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_188
timestamp 1626908933
transform 1 0 5472 0 -1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_41
timestamp 1626908933
transform 1 0 5520 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_241
timestamp 1626908933
transform 1 0 5520 0 1 333
box -32 -32 32 32
use L1M1_PR  L1M1_PR_50
timestamp 1626908933
transform 1 0 5520 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_52
timestamp 1626908933
transform 1 0 5424 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_270
timestamp 1626908933
transform 1 0 5520 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_272
timestamp 1626908933
transform 1 0 5424 0 1 333
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_0
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_12
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_62
timestamp 1626908933
transform 1 0 5760 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_181
timestamp 1626908933
transform 1 0 5760 0 1 0
box -38 -49 134 715
use M1M2_PR  M1M2_PR_17
timestamp 1626908933
transform 1 0 5808 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_217
timestamp 1626908933
transform 1 0 5808 0 1 555
box -32 -32 32 32
use L1M1_PR  L1M1_PR_19
timestamp 1626908933
transform 1 0 5712 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_239
timestamp 1626908933
transform 1 0 5712 0 1 555
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_61
timestamp 1626908933
transform 1 0 6624 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_180
timestamp 1626908933
transform 1 0 6624 0 1 0
box -38 -49 134 715
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_5
timestamp 1626908933
transform 1 0 6500 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_13
timestamp 1626908933
transform 1 0 6500 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_5
timestamp 1626908933
transform 1 0 6500 0 1 23
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_13
timestamp 1626908933
transform 1 0 6500 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_19
timestamp 1626908933
transform 1 0 6720 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_26
timestamp 1626908933
transform 1 0 5856 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_62
timestamp 1626908933
transform 1 0 6720 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_69
timestamp 1626908933
transform 1 0 5856 0 1 0
box -38 -49 806 715
use M1M2_PR  M1M2_PR_361
timestamp 1626908933
transform 1 0 7056 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_161
timestamp 1626908933
transform 1 0 7056 0 1 185
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_179
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_177
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_60
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_58
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_86
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_83
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_41
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_38
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_67
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_7
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_67
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_7
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_176
timestamp 1626908933
transform 1 0 8064 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_57
timestamp 1626908933
transform 1 0 8064 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_71
timestamp 1626908933
transform 1 0 7680 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_17
timestamp 1626908933
transform 1 0 7680 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_10
timestamp 1626908933
transform 1 0 8160 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_21
timestamp 1626908933
transform 1 0 8160 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_17
timestamp 1626908933
transform 1 0 7680 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_60
timestamp 1626908933
transform 1 0 7680 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_24
timestamp 1626908933
transform 1 0 5568 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_0
timestamp 1626908933
transform 1 0 5568 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_59
timestamp 1626908933
transform 1 0 8448 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_178
timestamp 1626908933
transform 1 0 8448 0 1 0
box -38 -49 134 715
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_4
timestamp 1626908933
transform 1 0 8900 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_12
timestamp 1626908933
transform 1 0 8900 0 1 16
box -100 -33 100 33
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_4
timestamp 1626908933
transform 1 0 8900 0 1 23
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_12
timestamp 1626908933
transform 1 0 8900 0 1 23
box -100 -26 100 26
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_8
timestamp 1626908933
transform 1 0 9024 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_9
timestamp 1626908933
transform 1 0 8928 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_51
timestamp 1626908933
transform 1 0 9024 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_52
timestamp 1626908933
transform 1 0 8928 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_12
timestamp 1626908933
transform 1 0 8640 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_13
timestamp 1626908933
transform 1 0 8544 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_66
timestamp 1626908933
transform 1 0 8640 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_67
timestamp 1626908933
transform 1 0 8544 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_40
timestamp 1626908933
transform 1 0 9696 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_85
timestamp 1626908933
transform 1 0 9696 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_20
timestamp 1626908933
transform 1 0 9792 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_24
timestamp 1626908933
transform 1 0 9792 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_81
timestamp 1626908933
transform 1 0 9792 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_85
timestamp 1626908933
transform 1 0 9792 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_65
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_70
timestamp 1626908933
transform 1 0 9984 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_184
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_189
timestamp 1626908933
transform 1 0 9984 0 -1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_359
timestamp 1626908933
transform 1 0 10032 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_159
timestamp 1626908933
transform 1 0 10032 0 1 185
box -32 -32 32 32
use L1M1_PR  L1M1_PR_344
timestamp 1626908933
transform 1 0 144 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_124
timestamp 1626908933
transform 1 0 144 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_380
timestamp 1626908933
transform 1 0 48 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_180
timestamp 1626908933
transform 1 0 48 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_381
timestamp 1626908933
transform 1 0 48 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_181
timestamp 1626908933
transform 1 0 48 0 1 1221
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_190
timestamp 1626908933
transform 1 0 192 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_71
timestamp 1626908933
transform 1 0 192 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_86
timestamp 1626908933
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_25
timestamp 1626908933
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_37
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_82
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_99
timestamp 1626908933
transform 1 0 336 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_299
timestamp 1626908933
transform 1 0 336 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_157
timestamp 1626908933
transform 1 0 528 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_377
timestamp 1626908933
transform 1 0 528 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_45
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_245
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_55
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_275
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_59
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_119
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_59
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_119
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use L1M1_PR  L1M1_PR_376
timestamp 1626908933
transform 1 0 2160 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_277
timestamp 1626908933
transform 1 0 2160 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_156
timestamp 1626908933
transform 1 0 2160 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_57
timestamp 1626908933
transform 1 0 2160 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_425
timestamp 1626908933
transform 1 0 2256 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_205
timestamp 1626908933
transform 1 0 2256 0 1 1073
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_191
timestamp 1626908933
transform 1 0 2304 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_72
timestamp 1626908933
transform 1 0 2304 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_276
timestamp 1626908933
transform 1 0 2448 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_56
timestamp 1626908933
transform 1 0 2448 0 1 1443
box -29 -23 29 23
use M1M2_PR  M1M2_PR_334
timestamp 1626908933
transform 1 0 2448 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_134
timestamp 1626908933
transform 1 0 2448 0 1 925
box -32 -32 32 32
use L1M1_PR  L1M1_PR_382
timestamp 1626908933
transform 1 0 2736 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_162
timestamp 1626908933
transform 1 0 2736 0 1 925
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_11
timestamp 1626908933
transform 1 0 2400 0 1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_23
timestamp 1626908933
transform 1 0 2400 0 1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_41
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_17
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_21
timestamp 1626908933
transform 1 0 2928 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_142
timestamp 1626908933
transform 1 0 3120 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_221
timestamp 1626908933
transform 1 0 2928 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_342
timestamp 1626908933
transform 1 0 3120 0 1 925
box -32 -32 32 32
use L1M1_PR  L1M1_PR_170
timestamp 1626908933
transform 1 0 3120 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_204
timestamp 1626908933
transform 1 0 2832 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_390
timestamp 1626908933
transform 1 0 3120 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_424
timestamp 1626908933
transform 1 0 2832 0 1 925
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_73
timestamp 1626908933
transform 1 0 3456 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_192
timestamp 1626908933
transform 1 0 3456 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_177
timestamp 1626908933
transform 1 0 3312 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_377
timestamp 1626908933
transform 1 0 3312 0 1 925
box -32 -32 32 32
use L1M1_PR  L1M1_PR_203
timestamp 1626908933
transform 1 0 3216 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_423
timestamp 1626908933
transform 1 0 3216 0 1 925
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_28
timestamp 1626908933
transform 1 0 3072 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_12
timestamp 1626908933
transform 1 0 3072 0 1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_53
timestamp 1626908933
transform 1 0 3792 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_253
timestamp 1626908933
transform 1 0 3792 0 1 1443
box -32 -32 32 32
use L1M1_PR  L1M1_PR_22
timestamp 1626908933
transform 1 0 3792 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_242
timestamp 1626908933
transform 1 0 3792 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_414
timestamp 1626908933
transform 1 0 3984 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_194
timestamp 1626908933
transform 1 0 3984 0 1 999
box -29 -23 29 23
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_112
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_52
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_112
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_52
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_193
timestamp 1626908933
transform 1 0 4224 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_74
timestamp 1626908933
transform 1 0 4224 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_87
timestamp 1626908933
transform 1 0 4032 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_26
timestamp 1626908933
transform 1 0 4032 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_14
timestamp 1626908933
transform 1 0 3552 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_3
timestamp 1626908933
transform 1 0 3552 0 1 1332
box -38 -49 518 715
use M1M2_PR  M1M2_PR_171
timestamp 1626908933
transform 1 0 4560 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_371
timestamp 1626908933
transform 1 0 4560 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_51
timestamp 1626908933
transform 1 0 4368 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_193
timestamp 1626908933
transform 1 0 4560 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_271
timestamp 1626908933
transform 1 0 4368 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_413
timestamp 1626908933
transform 1 0 4560 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_36
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_81
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_27
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_88
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_17
timestamp 1626908933
transform -1 0 4800 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_6
timestamp 1626908933
transform -1 0 4800 0 1 1332
box -38 -49 518 715
use M1M2_PR  M1M2_PR_40
timestamp 1626908933
transform 1 0 5520 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_43
timestamp 1626908933
transform 1 0 5136 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_240
timestamp 1626908933
transform 1 0 5520 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_243
timestamp 1626908933
transform 1 0 5136 0 1 777
box -32 -32 32 32
use L1M1_PR  L1M1_PR_53
timestamp 1626908933
transform 1 0 5136 0 1 777
box -29 -23 29 23
use L1M1_PR  L1M1_PR_273
timestamp 1626908933
transform 1 0 5136 0 1 777
box -29 -23 29 23
use L1M1_PR  L1M1_PR_66
timestamp 1626908933
transform 1 0 5136 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_286
timestamp 1626908933
transform 1 0 5136 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_9
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_21
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 710 715
use L1M1_PR  L1M1_PR_365
timestamp 1626908933
transform 1 0 5616 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_145
timestamp 1626908933
transform 1 0 5616 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_323
timestamp 1626908933
transform 1 0 5616 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_123
timestamp 1626908933
transform 1 0 5616 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_216
timestamp 1626908933
transform 1 0 5808 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_16
timestamp 1626908933
transform 1 0 5808 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_175
timestamp 1626908933
transform 1 0 5760 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_56
timestamp 1626908933
transform 1 0 5760 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_238
timestamp 1626908933
transform 1 0 6000 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_18
timestamp 1626908933
transform 1 0 6000 0 1 999
box -29 -23 29 23
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_105
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_45
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_105
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_45
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_78
timestamp 1626908933
transform 1 0 6624 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_17
timestamp 1626908933
transform 1 0 6624 0 1 1332
box -38 -49 230 715
use M1M2_PR  M1M2_PR_246
timestamp 1626908933
transform 1 0 6864 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_46
timestamp 1626908933
transform 1 0 6864 0 1 1221
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_174
timestamp 1626908933
transform 1 0 6816 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_55
timestamp 1626908933
transform 1 0 6816 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_18
timestamp 1626908933
transform 1 0 6912 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_25
timestamp 1626908933
transform 1 0 5856 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_61
timestamp 1626908933
transform 1 0 6912 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_68
timestamp 1626908933
transform 1 0 5856 0 1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_354
timestamp 1626908933
transform 1 0 8208 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_278
timestamp 1626908933
transform 1 0 7152 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_134
timestamp 1626908933
transform 1 0 8208 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_58
timestamp 1626908933
transform 1 0 7152 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_315
timestamp 1626908933
transform 1 0 7920 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_115
timestamp 1626908933
transform 1 0 7920 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_25
timestamp 1626908933
transform 1 0 7680 0 1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_1
timestamp 1626908933
transform 1 0 7680 0 1 1332
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_225
timestamp 1626908933
transform 1 0 8496 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_5
timestamp 1626908933
transform 1 0 8496 0 1 1221
box -29 -23 29 23
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_98
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_38
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_98
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_38
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use M1M2_PR  M1M2_PR_207
timestamp 1626908933
transform 1 0 9168 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_7
timestamp 1626908933
transform 1 0 9168 0 1 1221
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_194
timestamp 1626908933
transform 1 0 9600 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_75
timestamp 1626908933
transform 1 0 9600 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_89
timestamp 1626908933
transform 1 0 9792 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_28
timestamp 1626908933
transform 1 0 9792 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_80
timestamp 1626908933
transform 1 0 9696 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_35
timestamp 1626908933
transform 1 0 9696 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_195
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_76
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_382
timestamp 1626908933
transform 1 0 48 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_182
timestamp 1626908933
transform 1 0 48 0 1 2257
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_196
timestamp 1626908933
transform 1 0 192 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_77
timestamp 1626908933
transform 1 0 192 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_90
timestamp 1626908933
transform 1 0 0 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_29
timestamp 1626908933
transform 1 0 0 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_98
timestamp 1626908933
transform 1 0 336 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_298
timestamp 1626908933
transform 1 0 336 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_119
timestamp 1626908933
transform 1 0 432 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_339
timestamp 1626908933
transform 1 0 432 0 1 1665
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_30
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_90
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_30
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_90
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use L1M1_PR  L1M1_PR_9
timestamp 1626908933
transform 1 0 336 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_229
timestamp 1626908933
transform 1 0 336 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_381
timestamp 1626908933
transform 1 0 816 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_161
timestamp 1626908933
transform 1 0 816 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_384
timestamp 1626908933
transform 1 0 720 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_184
timestamp 1626908933
transform 1 0 720 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_133
timestamp 1626908933
transform 1 0 1104 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_333
timestamp 1626908933
transform 1 0 1104 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_132
timestamp 1626908933
transform 1 0 1104 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_332
timestamp 1626908933
transform 1 0 1104 0 1 2257
box -32 -32 32 32
use L1M1_PR  L1M1_PR_160
timestamp 1626908933
transform 1 0 1104 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_206
timestamp 1626908933
transform 1 0 1200 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_380
timestamp 1626908933
transform 1 0 1104 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_426
timestamp 1626908933
transform 1 0 1200 0 1 2257
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_30
timestamp 1626908933
transform 1 0 1344 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_91
timestamp 1626908933
transform 1 0 1344 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_5
timestamp 1626908933
transform 1 0 960 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_21
timestamp 1626908933
transform 1 0 960 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_8
timestamp 1626908933
transform -1 0 960 0 -1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_20
timestamp 1626908933
transform -1 0 960 0 -1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_16
timestamp 1626908933
transform 1 0 1536 0 -1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_5
timestamp 1626908933
transform 1 0 1536 0 -1 2664
box -38 -49 518 715
use M1M2_PR  M1M2_PR_44
timestamp 1626908933
transform 1 0 1872 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_244
timestamp 1626908933
transform 1 0 1872 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_24
timestamp 1626908933
transform 1 0 2016 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_8
timestamp 1626908933
transform 1 0 2016 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_34
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_79
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_78
timestamp 1626908933
transform 1 0 2400 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_197
timestamp 1626908933
transform 1 0 2400 0 -1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_54
timestamp 1626908933
transform 1 0 2448 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_274
timestamp 1626908933
transform 1 0 2448 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_25
timestamp 1626908933
transform 1 0 2736 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_245
timestamp 1626908933
transform 1 0 2736 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_29
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_5
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_20
timestamp 1626908933
transform 1 0 2928 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_220
timestamp 1626908933
transform 1 0 2928 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_23
timestamp 1626908933
transform 1 0 2832 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_243
timestamp 1626908933
transform 1 0 2832 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_24
timestamp 1626908933
transform 1 0 3696 0 1 1517
box -29 -23 29 23
use L1M1_PR  L1M1_PR_244
timestamp 1626908933
transform 1 0 3696 0 1 1517
box -29 -23 29 23
use L1M1_PR  L1M1_PR_196
timestamp 1626908933
transform 1 0 3888 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_416
timestamp 1626908933
transform 1 0 3888 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_147
timestamp 1626908933
transform 1 0 3120 0 1 1739
box -32 -32 32 32
use M1M2_PR  M1M2_PR_347
timestamp 1626908933
transform 1 0 3120 0 1 1739
box -32 -32 32 32
use L1M1_PR  L1M1_PR_21
timestamp 1626908933
transform 1 0 3024 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_241
timestamp 1626908933
transform 1 0 3024 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_174
timestamp 1626908933
transform 1 0 3216 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_207
timestamp 1626908933
transform 1 0 3312 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_394
timestamp 1626908933
transform 1 0 3216 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_427
timestamp 1626908933
transform 1 0 3312 0 1 1739
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_22
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_82
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_22
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_82
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use M1M2_PR  M1M2_PR_9
timestamp 1626908933
transform 1 0 3408 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_209
timestamp 1626908933
transform 1 0 3408 0 1 2109
box -32 -32 32 32
use L1M1_PR  L1M1_PR_412
timestamp 1626908933
transform 1 0 4560 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_249
timestamp 1626908933
transform 1 0 4656 0 1 1739
box -29 -23 29 23
use L1M1_PR  L1M1_PR_192
timestamp 1626908933
transform 1 0 4560 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_29
timestamp 1626908933
transform 1 0 4656 0 1 1739
box -29 -23 29 23
use M1M2_PR  M1M2_PR_370
timestamp 1626908933
transform 1 0 4560 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_170
timestamp 1626908933
transform 1 0 4560 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_285
timestamp 1626908933
transform 1 0 4368 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_65
timestamp 1626908933
transform 1 0 4368 0 1 2109
box -29 -23 29 23
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_6
timestamp 1626908933
transform -1 0 4992 0 -1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_14
timestamp 1626908933
transform -1 0 4992 0 -1 2664
box -38 -49 518 715
use L1M1_PR  L1M1_PR_247
timestamp 1626908933
transform 1 0 4752 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_27
timestamp 1626908933
transform 1 0 4752 0 1 2257
box -29 -23 29 23
use M1M2_PR  M1M2_PR_223
timestamp 1626908933
transform 1 0 4752 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_222
timestamp 1626908933
transform 1 0 4752 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_23
timestamp 1626908933
transform 1 0 4752 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_22
timestamp 1626908933
transform 1 0 4752 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_51
timestamp 1626908933
transform 1 0 5136 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_251
timestamp 1626908933
transform 1 0 5136 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_64
timestamp 1626908933
transform 1 0 5136 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_284
timestamp 1626908933
transform 1 0 5136 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_50
timestamp 1626908933
transform 1 0 5136 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_250
timestamp 1626908933
transform 1 0 5136 0 1 2109
box -32 -32 32 32
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_14
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_74
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_14
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_74
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_54
timestamp 1626908933
transform 1 0 4992 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_173
timestamp 1626908933
transform 1 0 4992 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_88
timestamp 1626908933
transform 1 0 5088 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_34
timestamp 1626908933
transform 1 0 5088 0 -1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_26
timestamp 1626908933
transform 1 0 5520 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_28
timestamp 1626908933
transform 1 0 5424 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_246
timestamp 1626908933
transform 1 0 5520 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_248
timestamp 1626908933
transform 1 0 5424 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_36
timestamp 1626908933
transform 1 0 5472 0 -1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_12
timestamp 1626908933
transform 1 0 5472 0 -1 2664
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_227
timestamp 1626908933
transform 1 0 5712 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_7
timestamp 1626908933
transform 1 0 5712 0 1 1591
box -29 -23 29 23
use M1M2_PR  M1M2_PR_219
timestamp 1626908933
transform 1 0 5808 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_19
timestamp 1626908933
transform 1 0 5808 0 1 1887
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_33
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_78
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_53
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_79
timestamp 1626908933
transform 1 0 7392 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_172
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_198
timestamp 1626908933
transform 1 0 7392 0 -1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_138
timestamp 1626908933
transform 1 0 7728 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_358
timestamp 1626908933
transform 1 0 7728 0 1 1665
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_6
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_66
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_6
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_66
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_16
timestamp 1626908933
transform 1 0 7680 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_70
timestamp 1626908933
transform 1 0 7680 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  sky130_fd_sc_hs__clkbuf_1_1
timestamp 1626908933
transform -1 0 8544 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  sky130_fd_sc_hs__clkbuf_1_0
timestamp 1626908933
transform -1 0 8544 0 -1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_226
timestamp 1626908933
transform 1 0 8112 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_6
timestamp 1626908933
transform 1 0 8112 0 1 1591
box -29 -23 29 23
use M1M2_PR  M1M2_PR_314
timestamp 1626908933
transform 1 0 7920 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_114
timestamp 1626908933
transform 1 0 7920 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_171
timestamp 1626908933
transform 1 0 8064 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_52
timestamp 1626908933
transform 1 0 8064 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_259
timestamp 1626908933
transform 1 0 8304 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_59
timestamp 1626908933
transform 1 0 8304 0 1 1887
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_170
timestamp 1626908933
transform 1 0 8544 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_51
timestamp 1626908933
transform 1 0 8544 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_65
timestamp 1626908933
transform 1 0 8640 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_11
timestamp 1626908933
transform 1 0 8640 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_50
timestamp 1626908933
transform 1 0 9024 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_7
timestamp 1626908933
transform 1 0 9024 0 -1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_292
timestamp 1626908933
transform 1 0 9264 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_72
timestamp 1626908933
transform 1 0 9264 0 1 1887
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_169
timestamp 1626908933
transform 1 0 9984 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_50
timestamp 1626908933
transform 1 0 9984 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_77
timestamp 1626908933
transform 1 0 9792 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_16
timestamp 1626908933
transform 1 0 9792 0 -1 2664
box -38 -49 230 715
use M1M2_PR  M1M2_PR_186
timestamp 1626908933
transform 1 0 240 0 1 2479
box -32 -32 32 32
use M1M2_PR  M1M2_PR_386
timestamp 1626908933
transform 1 0 240 0 1 2479
box -32 -32 32 32
use M1M2_PR  M1M2_PR_173
timestamp 1626908933
transform 1 0 144 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_185
timestamp 1626908933
transform 1 0 48 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_373
timestamp 1626908933
transform 1 0 144 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_385
timestamp 1626908933
transform 1 0 48 0 1 2775
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_31
timestamp 1626908933
transform 1 0 0 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_92
timestamp 1626908933
transform 1 0 0 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_80
timestamp 1626908933
transform 1 0 192 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_199
timestamp 1626908933
transform 1 0 192 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_251
timestamp 1626908933
transform 1 0 528 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_31
timestamp 1626908933
transform 1 0 528 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_225
timestamp 1626908933
transform 1 0 528 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_25
timestamp 1626908933
transform 1 0 528 0 1 2331
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_93
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_32
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_77
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_32
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_253
timestamp 1626908933
transform 1 0 624 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_33
timestamp 1626908933
transform 1 0 624 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_383
timestamp 1626908933
transform 1 0 720 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_224
timestamp 1626908933
transform 1 0 624 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_183
timestamp 1626908933
transform 1 0 720 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_24
timestamp 1626908933
transform 1 0 624 0 1 2923
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_200
timestamp 1626908933
transform 1 0 576 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_81
timestamp 1626908933
transform 1 0 576 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_69
timestamp 1626908933
transform 1 0 912 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_289
timestamp 1626908933
transform 1 0 912 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_57
timestamp 1626908933
transform 1 0 912 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_257
timestamp 1626908933
transform 1 0 912 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_71
timestamp 1626908933
transform 1 0 912 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_291
timestamp 1626908933
transform 1 0 912 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_30
timestamp 1626908933
transform 1 0 912 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_250
timestamp 1626908933
transform 1 0 912 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_200
timestamp 1626908933
transform 1 0 1104 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_420
timestamp 1626908933
transform 1 0 1104 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_4
timestamp 1626908933
transform 1 0 672 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_12
timestamp 1626908933
transform 1 0 672 0 1 2664
box -38 -49 518 715
use M1M2_PR  M1M2_PR_90
timestamp 1626908933
transform 1 0 1200 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_290
timestamp 1626908933
transform 1 0 1200 0 1 2997
box -32 -32 32 32
use L1M1_PR  L1M1_PR_115
timestamp 1626908933
transform 1 0 1200 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_335
timestamp 1626908933
transform 1 0 1200 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_55
timestamp 1626908933
transform 1 0 1392 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_255
timestamp 1626908933
transform 1 0 1392 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_32
timestamp 1626908933
transform 1 0 1968 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_199
timestamp 1626908933
transform 1 0 1872 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_252
timestamp 1626908933
transform 1 0 1968 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_419
timestamp 1626908933
transform 1 0 1872 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_208
timestamp 1626908933
transform 1 0 2256 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_428
timestamp 1626908933
transform 1 0 2256 0 1 2405
box -29 -23 29 23
use M1M2_PR  M1M2_PR_87
timestamp 1626908933
transform 1 0 2640 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_287
timestamp 1626908933
transform 1 0 2640 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_110
timestamp 1626908933
transform 1 0 2640 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_330
timestamp 1626908933
transform 1 0 2640 0 1 2331
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_58
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_118
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_58
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_118
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use M1M2_PR  M1M2_PR_139
timestamp 1626908933
transform 1 0 2160 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_339
timestamp 1626908933
transform 1 0 2160 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_166
timestamp 1626908933
transform 1 0 2160 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_386
timestamp 1626908933
transform 1 0 2160 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_167
timestamp 1626908933
transform 1 0 1584 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_387
timestamp 1626908933
transform 1 0 1584 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_138
timestamp 1626908933
transform 1 0 2160 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_338
timestamp 1626908933
transform 1 0 2160 0 1 2923
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_42
timestamp 1626908933
transform 1 0 1152 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_18
timestamp 1626908933
transform 1 0 1152 0 1 2664
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_146
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_346
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -32 -32 32 32
use L1M1_PR  L1M1_PR_175
timestamp 1626908933
transform 1 0 3024 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_395
timestamp 1626908933
transform 1 0 3024 0 1 2405
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_51
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_111
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_51
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_111
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use L1M1_PR  L1M1_PR_67
timestamp 1626908933
transform 1 0 2928 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_287
timestamp 1626908933
transform 1 0 2928 0 1 2775
box -29 -23 29 23
use M1M2_PR  M1M2_PR_80
timestamp 1626908933
transform 1 0 3216 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_280
timestamp 1626908933
transform 1 0 3216 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_8
timestamp 1626908933
transform 1 0 3408 0 1 2849
box -32 -32 32 32
use M1M2_PR  M1M2_PR_208
timestamp 1626908933
transform 1 0 3408 0 1 2849
box -32 -32 32 32
use M1M2_PR  M1M2_PR_52
timestamp 1626908933
transform 1 0 3792 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_252
timestamp 1626908933
transform 1 0 3792 0 1 2775
box -32 -32 32 32
use L1M1_PR  L1M1_PR_106
timestamp 1626908933
transform 1 0 3216 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_326
timestamp 1626908933
transform 1 0 3216 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_169
timestamp 1626908933
transform 1 0 4560 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_369
timestamp 1626908933
transform 1 0 4560 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_191
timestamp 1626908933
transform 1 0 4560 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_411
timestamp 1626908933
transform 1 0 4560 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_31
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_76
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_33
timestamp 1626908933
transform 1 0 5184 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_87
timestamp 1626908933
transform 1 0 5184 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_49
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_168
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_146
timestamp 1626908933
transform 1 0 5520 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_366
timestamp 1626908933
transform 1 0 5520 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_16  sky130_fd_sc_hs__clkbuf_16_0
timestamp 1626908933
transform 1 0 3072 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  sky130_fd_sc_hs__clkbuf_16_1
timestamp 1626908933
transform 1 0 3072 0 1 2664
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_122
timestamp 1626908933
transform 1 0 5616 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_322
timestamp 1626908933
transform 1 0 5616 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_18
timestamp 1626908933
transform 1 0 5808 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_218
timestamp 1626908933
transform 1 0 5808 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_20
timestamp 1626908933
transform 1 0 5904 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_240
timestamp 1626908933
transform 1 0 5904 0 1 2331
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_44
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_104
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_44
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_104
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use M1M2_PR  M1M2_PR_49
timestamp 1626908933
transform 1 0 6672 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_249
timestamp 1626908933
transform 1 0 6672 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_121
timestamp 1626908933
transform 1 0 5616 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_321
timestamp 1626908933
transform 1 0 5616 0 1 2997
box -32 -32 32 32
use L1M1_PR  L1M1_PR_8
timestamp 1626908933
transform 1 0 6000 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_228
timestamp 1626908933
transform 1 0 6000 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_144
timestamp 1626908933
transform 1 0 5616 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_364
timestamp 1626908933
transform 1 0 5616 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_104
timestamp 1626908933
transform 1 0 7632 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_304
timestamp 1626908933
transform 1 0 7632 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_60
timestamp 1626908933
transform 1 0 7056 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_126
timestamp 1626908933
transform 1 0 8208 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_280
timestamp 1626908933
transform 1 0 7056 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_346
timestamp 1626908933
transform 1 0 8208 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_307
timestamp 1626908933
transform 1 0 7536 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_87
timestamp 1626908933
transform 1 0 7536 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_294
timestamp 1626908933
transform 1 0 8208 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_74
timestamp 1626908933
transform 1 0 8208 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_295
timestamp 1626908933
transform 1 0 7344 0 1 2849
box -29 -23 29 23
use L1M1_PR  L1M1_PR_75
timestamp 1626908933
transform 1 0 7344 0 1 2849
box -29 -23 29 23
use M2M3_PR  M2M3_PR_11
timestamp 1626908933
transform 1 0 7920 0 1 2965
box -33 -37 33 37
use M2M3_PR  M2M3_PR_5
timestamp 1626908933
transform 1 0 7920 0 1 2965
box -33 -37 33 37
use M1M2_PR  M1M2_PR_267
timestamp 1626908933
transform 1 0 8112 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_67
timestamp 1626908933
transform 1 0 8112 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_305
timestamp 1626908933
transform 1 0 7536 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_85
timestamp 1626908933
transform 1 0 7536 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_303
timestamp 1626908933
transform 1 0 7632 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_103
timestamp 1626908933
transform 1 0 7632 0 1 2997
box -32 -32 32 32
use L1M1_PR  L1M1_PR_347
timestamp 1626908933
transform 1 0 7824 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_127
timestamp 1626908933
transform 1 0 7824 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_356
timestamp 1626908933
transform 1 0 7920 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_136
timestamp 1626908933
transform 1 0 7920 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_313
timestamp 1626908933
transform 1 0 7920 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_113
timestamp 1626908933
transform 1 0 7920 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_4
timestamp 1626908933
transform 1 0 7488 0 1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_7
timestamp 1626908933
transform 1 0 8160 0 1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_16
timestamp 1626908933
transform 1 0 7488 0 1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_19
timestamp 1626908933
transform 1 0 8160 0 1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_37
timestamp 1626908933
transform 1 0 5568 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_13
timestamp 1626908933
transform 1 0 5568 0 1 2664
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_351
timestamp 1626908933
transform 1 0 8496 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_131
timestamp 1626908933
transform 1 0 8496 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_307
timestamp 1626908933
transform 1 0 8688 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_107
timestamp 1626908933
transform 1 0 8688 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_302
timestamp 1626908933
transform 1 0 8496 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_102
timestamp 1626908933
transform 1 0 8496 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_293
timestamp 1626908933
transform 1 0 8304 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_73
timestamp 1626908933
transform 1 0 8304 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_258
timestamp 1626908933
transform 1 0 8304 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_58
timestamp 1626908933
transform 1 0 8304 0 1 2997
box -32 -32 32 32
use L1M1_PR  L1M1_PR_345
timestamp 1626908933
transform 1 0 8496 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_125
timestamp 1626908933
transform 1 0 8496 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_301
timestamp 1626908933
transform 1 0 8496 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_101
timestamp 1626908933
transform 1 0 8496 0 1 2997
box -32 -32 32 32
use M2M3_PR  M2M3_PR_10
timestamp 1626908933
transform 1 0 8592 0 1 2965
box -33 -37 33 37
use M2M3_PR  M2M3_PR_4
timestamp 1626908933
transform 1 0 8592 0 1 2965
box -33 -37 33 37
use L1M1_PR  L1M1_PR_353
timestamp 1626908933
transform 1 0 8592 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_133
timestamp 1626908933
transform 1 0 8592 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_310
timestamp 1626908933
transform 1 0 8592 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_110
timestamp 1626908933
transform 1 0 8592 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_48
timestamp 1626908933
transform 1 0 8832 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_167
timestamp 1626908933
transform 1 0 8832 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_183
timestamp 1626908933
transform 1 0 8784 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_403
timestamp 1626908933
transform 1 0 8784 0 1 2997
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_37
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_97
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_37
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_97
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_6
timestamp 1626908933
transform 1 0 8928 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_49
timestamp 1626908933
transform 1 0 8928 0 1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_357
timestamp 1626908933
transform 1 0 9456 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_157
timestamp 1626908933
transform 1 0 9456 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_201
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_82
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_94
timestamp 1626908933
transform 1 0 9792 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_33
timestamp 1626908933
transform 1 0 9792 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_75
timestamp 1626908933
transform 1 0 9696 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_30
timestamp 1626908933
transform 1 0 9696 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_83
timestamp 1626908933
transform 1 0 0 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_202
timestamp 1626908933
transform 1 0 0 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_123
timestamp 1626908933
transform 1 0 144 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_343
timestamp 1626908933
transform 1 0 144 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_97
timestamp 1626908933
transform 1 0 336 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_297
timestamp 1626908933
transform 1 0 336 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_159
timestamp 1626908933
transform 1 0 528 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_379
timestamp 1626908933
transform 1 0 528 0 1 3663
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_29
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_89
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_29
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_89
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_54
timestamp 1626908933
transform 1 0 1392 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_254
timestamp 1626908933
transform 1 0 1392 0 1 3441
box -32 -32 32 32
use L1M1_PR  L1M1_PR_68
timestamp 1626908933
transform 1 0 1680 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_288
timestamp 1626908933
transform 1 0 1680 0 1 3441
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_20
timestamp 1626908933
transform 1 0 2016 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_4
timestamp 1626908933
transform 1 0 2016 0 -1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_158
timestamp 1626908933
transform 1 0 2160 0 1 3589
box -29 -23 29 23
use L1M1_PR  L1M1_PR_209
timestamp 1626908933
transform 1 0 2256 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_378
timestamp 1626908933
transform 1 0 2160 0 1 3589
box -29 -23 29 23
use L1M1_PR  L1M1_PR_429
timestamp 1626908933
transform 1 0 2256 0 1 3737
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_29
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_74
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_43
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_97
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_84
timestamp 1626908933
transform 1 0 2400 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_203
timestamp 1626908933
transform 1 0 2400 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_30
timestamp 1626908933
transform 1 0 96 0 -1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_6
timestamp 1626908933
transform 1 0 96 0 -1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_34
timestamp 1626908933
transform 1 0 2976 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_95
timestamp 1626908933
transform 1 0 2976 0 -1 3996
box -38 -49 230 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_21
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_81
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_21
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_81
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_79
timestamp 1626908933
transform 1 0 3216 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_279
timestamp 1626908933
transform 1 0 3216 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_105
timestamp 1626908933
transform 1 0 3216 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_325
timestamp 1626908933
transform 1 0 3216 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_168
timestamp 1626908933
transform 1 0 4560 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_368
timestamp 1626908933
transform 1 0 4560 0 1 3071
box -32 -32 32 32
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_13
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_73
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_13
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_73
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_1
timestamp 1626908933
transform 1 0 5040 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_201
timestamp 1626908933
transform 1 0 5040 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3
timestamp 1626908933
transform 1 0 4752 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_203
timestamp 1626908933
transform 1 0 4752 0 1 3737
box -32 -32 32 32
use L1M1_PR  L1M1_PR_132
timestamp 1626908933
transform 1 0 5424 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_352
timestamp 1626908933
transform 1 0 5424 0 1 3663
box -29 -23 29 23
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_2
timestamp 1626908933
transform -1 0 5856 0 -1 3996
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_0
timestamp 1626908933
transform -1 0 5856 0 -1 3996
box -38 -49 2726 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_35
timestamp 1626908933
transform 1 0 5856 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_96
timestamp 1626908933
transform 1 0 5856 0 -1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1
timestamp 1626908933
transform 1 0 5808 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_221
timestamp 1626908933
transform 1 0 5808 0 1 3737
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_85
timestamp 1626908933
transform 1 0 6048 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_204
timestamp 1626908933
transform 1 0 6048 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_63
timestamp 1626908933
transform 1 0 6096 0 1 3515
box -29 -23 29 23
use L1M1_PR  L1M1_PR_283
timestamp 1626908933
transform 1 0 6096 0 1 3515
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_10
timestamp 1626908933
transform -1 0 6816 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_22
timestamp 1626908933
transform -1 0 6816 0 -1 3996
box -38 -49 710 715
use M1M2_PR  M1M2_PR_309
timestamp 1626908933
transform 1 0 6288 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_109
timestamp 1626908933
transform 1 0 6288 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_248
timestamp 1626908933
transform 1 0 6672 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_48
timestamp 1626908933
transform 1 0 6672 0 1 3515
box -32 -32 32 32
use L1M1_PR  L1M1_PR_405
timestamp 1626908933
transform 1 0 6864 0 1 3515
box -29 -23 29 23
use L1M1_PR  L1M1_PR_185
timestamp 1626908933
transform 1 0 6864 0 1 3515
box -29 -23 29 23
use L1M1_PR  L1M1_PR_361
timestamp 1626908933
transform 1 0 6384 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_141
timestamp 1626908933
transform 1 0 6384 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_308
timestamp 1626908933
transform 1 0 6288 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_108
timestamp 1626908933
transform 1 0 6288 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_349
timestamp 1626908933
transform 1 0 6480 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_129
timestamp 1626908933
transform 1 0 6480 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_279
timestamp 1626908933
transform 1 0 6768 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_59
timestamp 1626908933
transform 1 0 6768 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_247
timestamp 1626908933
transform 1 0 6768 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_47
timestamp 1626908933
transform 1 0 6768 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_317
timestamp 1626908933
transform 1 0 6384 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_117
timestamp 1626908933
transform 1 0 6384 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_1
timestamp 1626908933
transform -1 0 7488 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_13
timestamp 1626908933
transform -1 0 7488 0 -1 3996
box -38 -49 710 715
use M1M2_PR  M1M2_PR_360
timestamp 1626908933
transform 1 0 7056 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_160
timestamp 1626908933
transform 1 0 7056 0 1 3515
box -32 -32 32 32
use L1M1_PR  L1M1_PR_359
timestamp 1626908933
transform 1 0 7056 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_348
timestamp 1626908933
transform 1 0 7152 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_139
timestamp 1626908933
transform 1 0 7056 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_128
timestamp 1626908933
transform 1 0 7152 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_316
timestamp 1626908933
transform 1 0 7056 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_116
timestamp 1626908933
transform 1 0 7056 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_305
timestamp 1626908933
transform 1 0 7248 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_105
timestamp 1626908933
transform 1 0 7248 0 1 3663
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_65
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_5
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_65
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_5
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_317
timestamp 1626908933
transform 1 0 7440 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_97
timestamp 1626908933
transform 1 0 7440 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_325
timestamp 1626908933
transform 1 0 7728 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_275
timestamp 1626908933
transform 1 0 7536 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_125
timestamp 1626908933
transform 1 0 7728 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_75
timestamp 1626908933
transform 1 0 7536 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_73
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_28
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_3
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_1
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 614 715
use M1M2_PR  M1M2_PR_112
timestamp 1626908933
transform 1 0 7920 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_312
timestamp 1626908933
transform 1 0 7920 0 1 3589
box -32 -32 32 32
use L1M1_PR  L1M1_PR_135
timestamp 1626908933
transform 1 0 7920 0 1 3589
box -29 -23 29 23
use L1M1_PR  L1M1_PR_148
timestamp 1626908933
transform 1 0 8016 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_355
timestamp 1626908933
transform 1 0 7920 0 1 3589
box -29 -23 29 23
use L1M1_PR  L1M1_PR_368
timestamp 1626908933
transform 1 0 8016 0 1 3737
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_36
timestamp 1626908933
transform 1 0 8160 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_97
timestamp 1626908933
transform 1 0 8160 0 -1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_184
timestamp 1626908933
transform 1 0 8112 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_404
timestamp 1626908933
transform 1 0 8112 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_269
timestamp 1626908933
transform 1 0 8400 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_69
timestamp 1626908933
transform 1 0 8400 0 1 3071
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_205
timestamp 1626908933
transform 1 0 8352 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_86
timestamp 1626908933
transform 1 0 8352 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_367
timestamp 1626908933
transform 1 0 8592 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_350
timestamp 1626908933
transform 1 0 8592 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_147
timestamp 1626908933
transform 1 0 8592 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_130
timestamp 1626908933
transform 1 0 8592 0 1 3441
box -29 -23 29 23
use M1M2_PR  M1M2_PR_306
timestamp 1626908933
transform 1 0 8688 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_106
timestamp 1626908933
transform 1 0 8688 0 1 3441
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_47
timestamp 1626908933
transform 1 0 9120 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_166
timestamp 1626908933
transform 1 0 9120 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__clkinv_4  sky130_fd_sc_hs__clkinv_4_0
timestamp 1626908933
transform 1 0 8448 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__clkinv_4  sky130_fd_sc_hs__clkinv_4_1
timestamp 1626908933
transform 1 0 8448 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_165
timestamp 1626908933
transform 1 0 9984 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_46
timestamp 1626908933
transform 1 0 9984 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_43
timestamp 1626908933
transform 1 0 9216 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_0
timestamp 1626908933
transform 1 0 9216 0 -1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_358
timestamp 1626908933
transform 1 0 10032 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_158
timestamp 1626908933
transform 1 0 10032 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_388
timestamp 1626908933
transform 1 0 48 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_387
timestamp 1626908933
transform 1 0 48 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_188
timestamp 1626908933
transform 1 0 48 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_187
timestamp 1626908933
transform 1 0 48 0 1 3885
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_206
timestamp 1626908933
transform 1 0 192 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_87
timestamp 1626908933
transform 1 0 192 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_389
timestamp 1626908933
transform 1 0 240 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_296
timestamp 1626908933
transform 1 0 336 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_189
timestamp 1626908933
transform 1 0 240 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_96
timestamp 1626908933
transform 1 0 336 0 1 4403
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_207
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_88
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_72
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_27
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_98
timestamp 1626908933
transform 1 0 0 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_37
timestamp 1626908933
transform 1 0 0 0 1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_129
timestamp 1626908933
transform 1 0 720 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_329
timestamp 1626908933
transform 1 0 720 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_152
timestamp 1626908933
transform 1 0 624 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_210
timestamp 1626908933
transform 1 0 720 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_372
timestamp 1626908933
transform 1 0 624 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_430
timestamp 1626908933
transform 1 0 720 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_17
timestamp 1626908933
transform 1 0 480 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_1
timestamp 1626908933
transform 1 0 480 0 1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_374
timestamp 1626908933
transform 1 0 1008 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_154
timestamp 1626908933
transform 1 0 1008 0 1 4107
box -29 -23 29 23
use M1M2_PR  M1M2_PR_331
timestamp 1626908933
transform 1 0 1008 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_131
timestamp 1626908933
transform 1 0 1008 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_431
timestamp 1626908933
transform 1 0 1104 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_211
timestamp 1626908933
transform 1 0 1104 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_289
timestamp 1626908933
transform 1 0 1200 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_89
timestamp 1626908933
transform 1 0 1200 0 1 4403
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_208
timestamp 1626908933
transform 1 0 1248 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_89
timestamp 1626908933
transform 1 0 1248 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_114
timestamp 1626908933
transform 1 0 1680 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_334
timestamp 1626908933
transform 1 0 1680 0 1 4403
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_57
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_117
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_57
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_117
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_18
timestamp 1626908933
transform 1 0 864 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_2
timestamp 1626908933
transform 1 0 1344 0 1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_2
timestamp 1626908933
transform 1 0 864 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_0
timestamp 1626908933
transform 1 0 1344 0 1 3996
box -38 -49 614 715
use L1M1_PR  L1M1_PR_327
timestamp 1626908933
transform 1 0 1776 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_107
timestamp 1626908933
transform 1 0 1776 0 1 4255
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_164
timestamp 1626908933
transform 1 0 1920 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_45
timestamp 1626908933
transform 1 0 1920 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_81
timestamp 1626908933
transform 1 0 2016 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_38
timestamp 1626908933
transform 1 0 2016 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_286
timestamp 1626908933
transform 1 0 2640 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_86
timestamp 1626908933
transform 1 0 2640 0 1 4403
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_44
timestamp 1626908933
transform 1 0 2784 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_163
timestamp 1626908933
transform 1 0 2784 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_81
timestamp 1626908933
transform 1 0 3024 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_281
timestamp 1626908933
transform 1 0 3024 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_27
timestamp 1626908933
transform 1 0 3312 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_227
timestamp 1626908933
transform 1 0 3312 0 1 4403
box -32 -32 32 32
use L1M1_PR  L1M1_PR_34
timestamp 1626908933
transform 1 0 3504 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_254
timestamp 1626908933
transform 1 0 3504 0 1 4403
box -29 -23 29 23
use M2M3_PR  M2M3_PR_3
timestamp 1626908933
transform 1 0 3216 0 1 4185
box -33 -37 33 37
use M2M3_PR  M2M3_PR_9
timestamp 1626908933
transform 1 0 3216 0 1 4185
box -33 -37 33 37
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_9
timestamp 1626908933
transform 1 0 3264 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_1
timestamp 1626908933
transform 1 0 3264 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_41
timestamp 1626908933
transform 1 0 2880 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_95
timestamp 1626908933
transform 1 0 2880 0 1 3996
box -38 -49 422 715
use M2M3_PR  M2M3_PR_2
timestamp 1626908933
transform 1 0 3888 0 1 4185
box -33 -37 33 37
use M2M3_PR  M2M3_PR_8
timestamp 1626908933
transform 1 0 3888 0 1 4185
box -33 -37 33 37
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_50
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_110
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_50
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_110
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_78
timestamp 1626908933
transform 1 0 3888 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_278
timestamp 1626908933
transform 1 0 3888 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_104
timestamp 1626908933
transform 1 0 4272 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_197
timestamp 1626908933
transform 1 0 3792 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_324
timestamp 1626908933
transform 1 0 4272 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_417
timestamp 1626908933
transform 1 0 3792 0 1 4477
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_19
timestamp 1626908933
transform -1 0 4608 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_8
timestamp 1626908933
transform -1 0 4608 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_0
timestamp 1626908933
transform 1 0 3744 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_2
timestamp 1626908933
transform 1 0 3744 0 1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_2
timestamp 1626908933
transform 1 0 4752 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_167
timestamp 1626908933
transform 1 0 4560 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_202
timestamp 1626908933
transform 1 0 4752 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_367
timestamp 1626908933
transform 1 0 4560 0 1 4477
box -32 -32 32 32
use L1M1_PR  L1M1_PR_2
timestamp 1626908933
transform 1 0 4464 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_222
timestamp 1626908933
transform 1 0 4464 0 1 4107
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_26
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_71
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_43
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_162
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_32
timestamp 1626908933
transform 1 0 5184 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_75
timestamp 1626908933
transform 1 0 5184 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_35
timestamp 1626908933
transform 1 0 4608 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_89
timestamp 1626908933
transform 1 0 4608 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_15
timestamp 1626908933
transform 1 0 5952 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_76
timestamp 1626908933
transform 1 0 5952 0 1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_402
timestamp 1626908933
transform 1 0 6192 0 1 3811
box -29 -23 29 23
use L1M1_PR  L1M1_PR_282
timestamp 1626908933
transform 1 0 6096 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_182
timestamp 1626908933
transform 1 0 6192 0 1 3811
box -29 -23 29 23
use L1M1_PR  L1M1_PR_62
timestamp 1626908933
transform 1 0 6096 0 1 3885
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_161
timestamp 1626908933
transform 1 0 6144 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_42
timestamp 1626908933
transform 1 0 6144 0 1 3996
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_103
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_43
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_103
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_43
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_83
timestamp 1626908933
transform 1 0 6240 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_29
timestamp 1626908933
transform 1 0 6240 0 1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_61
timestamp 1626908933
transform 1 0 6768 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_281
timestamp 1626908933
transform 1 0 6768 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_369
timestamp 1626908933
transform 1 0 6960 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_318
timestamp 1626908933
transform 1 0 7440 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_149
timestamp 1626908933
transform 1 0 6960 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_98
timestamp 1626908933
transform 1 0 7440 0 1 3885
box -29 -23 29 23
use M1M2_PR  M1M2_PR_324
timestamp 1626908933
transform 1 0 7728 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_277
timestamp 1626908933
transform 1 0 7344 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_124
timestamp 1626908933
transform 1 0 7728 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_77
timestamp 1626908933
transform 1 0 7344 0 1 3885
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_3
timestamp 1626908933
transform -1 0 9312 0 1 3996
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_1
timestamp 1626908933
transform -1 0 9312 0 1 3996
box -38 -49 2726 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_36
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_96
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_36
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_96
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_6
timestamp 1626908933
transform 1 0 9168 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_206
timestamp 1626908933
transform 1 0 9168 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_5
timestamp 1626908933
transform 1 0 8784 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_205
timestamp 1626908933
transform 1 0 8784 0 1 4403
box -32 -32 32 32
use L1M1_PR  L1M1_PR_219
timestamp 1626908933
transform 1 0 8880 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_439
timestamp 1626908933
transform 1 0 8880 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_224
timestamp 1626908933
transform 1 0 9264 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_4
timestamp 1626908933
transform 1 0 9264 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_356
timestamp 1626908933
transform 1 0 9456 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_156
timestamp 1626908933
transform 1 0 9456 0 1 4477
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_55
timestamp 1626908933
transform 1 0 9312 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1
timestamp 1626908933
transform 1 0 9312 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_25
timestamp 1626908933
transform 1 0 9696 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_70
timestamp 1626908933
transform 1 0 9696 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_154
timestamp 1626908933
transform 1 0 9744 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_199
timestamp 1626908933
transform 1 0 9840 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_354
timestamp 1626908933
transform 1 0 9744 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_399
timestamp 1626908933
transform 1 0 9840 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_90
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_209
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_155
timestamp 1626908933
transform 1 0 10032 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_355
timestamp 1626908933
transform 1 0 10032 0 1 4477
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_38
timestamp 1626908933
transform 1 0 9792 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_99
timestamp 1626908933
transform 1 0 9792 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_41
timestamp 1626908933
transform 1 0 0 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_102
timestamp 1626908933
transform 1 0 0 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_91
timestamp 1626908933
transform 1 0 0 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_94
timestamp 1626908933
transform 1 0 192 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_210
timestamp 1626908933
transform 1 0 0 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_213
timestamp 1626908933
transform 1 0 192 0 1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_122
timestamp 1626908933
transform 1 0 144 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_342
timestamp 1626908933
transform 1 0 144 0 1 4995
box -29 -23 29 23
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_88
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_28
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_88
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_28
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_373
timestamp 1626908933
transform 1 0 528 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_153
timestamp 1626908933
transform 1 0 528 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_295
timestamp 1626908933
transform 1 0 336 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_95
timestamp 1626908933
transform 1 0 336 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_67
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_22
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_128
timestamp 1626908933
transform 1 0 720 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_328
timestamp 1626908933
transform 1 0 720 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_56
timestamp 1626908933
transform 1 0 912 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_256
timestamp 1626908933
transform 1 0 912 0 1 4773
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_116
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_56
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_116
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_56
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use L1M1_PR  L1M1_PR_290
timestamp 1626908933
transform 1 0 1680 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_70
timestamp 1626908933
transform 1 0 1680 0 1 4773
box -29 -23 29 23
use M1M2_PR  M1M2_PR_263
timestamp 1626908933
transform 1 0 1872 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_63
timestamp 1626908933
transform 1 0 1872 0 1 5217
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_160
timestamp 1626908933
transform 1 0 2016 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_41
timestamp 1626908933
transform 1 0 2016 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_261
timestamp 1626908933
transform 1 0 2160 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_61
timestamp 1626908933
transform 1 0 2160 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_298
timestamp 1626908933
transform 1 0 2640 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_296
timestamp 1626908933
transform 1 0 2640 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_78
timestamp 1626908933
transform 1 0 2640 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_76
timestamp 1626908933
transform 1 0 2640 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_69
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_24
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_100
timestamp 1626908933
transform 1 0 2112 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_46
timestamp 1626908933
transform 1 0 2112 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_6
timestamp 1626908933
transform 1 0 2592 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_18
timestamp 1626908933
transform 1 0 2592 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_43
timestamp 1626908933
transform 1 0 96 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_32
timestamp 1626908933
transform 1 0 2304 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_31
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_19
timestamp 1626908933
transform 1 0 96 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_8
timestamp 1626908933
transform 1 0 2304 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_7
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_35
timestamp 1626908933
transform 1 0 3024 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_37
timestamp 1626908933
transform 1 0 2928 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_255
timestamp 1626908933
transform 1 0 3024 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_257
timestamp 1626908933
transform 1 0 2928 0 1 4995
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_20
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_80
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_20
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_80
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_39
timestamp 1626908933
transform 1 0 3264 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_100
timestamp 1626908933
transform 1 0 3264 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_92
timestamp 1626908933
transform 1 0 3456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_211
timestamp 1626908933
transform 1 0 3456 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_26
timestamp 1626908933
transform 1 0 3312 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_226
timestamp 1626908933
transform 1 0 3312 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_11
timestamp 1626908933
transform 1 0 3216 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_231
timestamp 1626908933
transform 1 0 3216 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_15
timestamp 1626908933
transform 1 0 3552 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_4
timestamp 1626908933
transform 1 0 3552 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_40
timestamp 1626908933
transform 1 0 4032 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_101
timestamp 1626908933
transform 1 0 4032 0 -1 5328
box -38 -49 230 715
use M1M2_PR  M1M2_PR_175
timestamp 1626908933
transform 1 0 3792 0 1 4921
box -32 -32 32 32
use M1M2_PR  M1M2_PR_375
timestamp 1626908933
transform 1 0 3792 0 1 4921
box -32 -32 32 32
use L1M1_PR  L1M1_PR_36
timestamp 1626908933
transform 1 0 3696 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_195
timestamp 1626908933
transform 1 0 3888 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_256
timestamp 1626908933
transform 1 0 3696 0 1 4921
box -29 -23 29 23
use L1M1_PR  L1M1_PR_415
timestamp 1626908933
transform 1 0 3888 0 1 4995
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_49
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_109
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_49
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_109
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_8
timestamp 1626908933
transform 1 0 4224 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_0
timestamp 1626908933
transform 1 0 4224 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_34
timestamp 1626908933
transform 1 0 4224 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_77
timestamp 1626908933
transform 1 0 4224 0 1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_166
timestamp 1626908933
transform 1 0 4560 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_366
timestamp 1626908933
transform 1 0 4560 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_39
timestamp 1626908933
transform 1 0 4464 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_190
timestamp 1626908933
transform 1 0 4656 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_202
timestamp 1626908933
transform 1 0 4848 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_259
timestamp 1626908933
transform 1 0 4464 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_410
timestamp 1626908933
transform 1 0 4656 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_422
timestamp 1626908933
transform 1 0 4848 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_220
timestamp 1626908933
transform 1 0 5040 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_0
timestamp 1626908933
transform 1 0 5040 0 1 4773
box -29 -23 29 23
use M1M2_PR  M1M2_PR_200
timestamp 1626908933
transform 1 0 5040 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_0
timestamp 1626908933
transform 1 0 5040 0 1 4773
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_66
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_21
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_72
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_12
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_72
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_12
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_20
timestamp 1626908933
transform -1 0 5184 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_9
timestamp 1626908933
transform -1 0 5184 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_31
timestamp 1626908933
transform 1 0 5184 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_74
timestamp 1626908933
transform 1 0 5184 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_5
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_17
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 710 715
use M1M2_PR  M1M2_PR_229
timestamp 1626908933
transform 1 0 5328 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_29
timestamp 1626908933
transform 1 0 5328 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_28
timestamp 1626908933
transform 1 0 6048 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_82
timestamp 1626908933
transform 1 0 6048 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_40
timestamp 1626908933
transform 1 0 5952 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_159
timestamp 1626908933
transform 1 0 5952 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_11
timestamp 1626908933
transform 1 0 6192 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_211
timestamp 1626908933
transform 1 0 6192 0 1 5217
box -32 -32 32 32
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_42
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_102
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_42
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_102
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_24
timestamp 1626908933
transform 1 0 6432 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_67
timestamp 1626908933
transform 1 0 6432 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_23
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_68
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_14
timestamp 1626908933
transform 1 0 7200 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_75
timestamp 1626908933
transform 1 0 7200 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_38
timestamp 1626908933
transform 1 0 7584 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_39
timestamp 1626908933
transform 1 0 7392 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_157
timestamp 1626908933
transform 1 0 7584 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_158
timestamp 1626908933
transform 1 0 7392 0 -1 5328
box -38 -49 134 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_4
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_64
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_4
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_64
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_16
timestamp 1626908933
transform 1 0 7680 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_59
timestamp 1626908933
transform 1 0 7680 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_38
timestamp 1626908933
transform 1 0 7680 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_26
timestamp 1626908933
transform 1 0 5760 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_14
timestamp 1626908933
transform 1 0 7680 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_2
timestamp 1626908933
transform 1 0 5760 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_74
timestamp 1626908933
transform 1 0 8448 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_13
timestamp 1626908933
transform 1 0 8448 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_64
timestamp 1626908933
transform 1 0 8640 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_10
timestamp 1626908933
transform 1 0 8640 0 -1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_4
timestamp 1626908933
transform 1 0 8784 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_204
timestamp 1626908933
transform 1 0 8784 0 1 4773
box -32 -32 32 32
use L1M1_PR  L1M1_PR_3
timestamp 1626908933
transform 1 0 9072 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_223
timestamp 1626908933
transform 1 0 9072 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_201
timestamp 1626908933
transform 1 0 9072 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_421
timestamp 1626908933
transform 1 0 9072 0 1 4995
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_35
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_95
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_35
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_95
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__clkinv_2  sky130_fd_sc_hs__clkinv_2_1
timestamp 1626908933
transform 1 0 9024 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__clkinv_2  sky130_fd_sc_hs__clkinv_2_0
timestamp 1626908933
transform 1 0 9024 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_214
timestamp 1626908933
transform 1 0 9600 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_156
timestamp 1626908933
transform 1 0 9408 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_95
timestamp 1626908933
transform 1 0 9600 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_37
timestamp 1626908933
transform 1 0 9408 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_54
timestamp 1626908933
transform 1 0 9504 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_0
timestamp 1626908933
transform 1 0 9504 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_20
timestamp 1626908933
transform 1 0 9696 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_65
timestamp 1626908933
transform 1 0 9696 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_36
timestamp 1626908933
transform 1 0 9888 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_155
timestamp 1626908933
transform 1 0 9888 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_93
timestamp 1626908933
transform 1 0 9984 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_96
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_212
timestamp 1626908933
transform 1 0 9984 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_215
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_42
timestamp 1626908933
transform 1 0 9792 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_103
timestamp 1626908933
transform 1 0 9792 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_97
timestamp 1626908933
transform 1 0 0 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_216
timestamp 1626908933
transform 1 0 0 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_94
timestamp 1626908933
transform 1 0 336 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_294
timestamp 1626908933
transform 1 0 336 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_118
timestamp 1626908933
transform 1 0 432 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_338
timestamp 1626908933
transform 1 0 432 0 1 5661
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_27
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_87
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_27
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_87
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_155
timestamp 1626908933
transform 1 0 816 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_375
timestamp 1626908933
transform 1 0 816 0 1 5587
box -29 -23 29 23
use M1M2_PR  M1M2_PR_130
timestamp 1626908933
transform 1 0 1008 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_330
timestamp 1626908933
transform 1 0 1008 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_45
timestamp 1626908933
transform 1 0 2112 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_99
timestamp 1626908933
transform 1 0 2112 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_35
timestamp 1626908933
transform 1 0 2016 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_154
timestamp 1626908933
transform 1 0 2016 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_60
timestamp 1626908933
transform 1 0 2160 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_260
timestamp 1626908933
transform 1 0 2160 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_77
timestamp 1626908933
transform 1 0 2160 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_297
timestamp 1626908933
transform 1 0 2160 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_333
timestamp 1626908933
transform 1 0 2352 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_113
timestamp 1626908933
transform 1 0 2352 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_64
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_19
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_397
timestamp 1626908933
transform 1 0 2736 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_177
timestamp 1626908933
transform 1 0 2736 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_285
timestamp 1626908933
transform 1 0 2640 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_85
timestamp 1626908933
transform 1 0 2640 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_217
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_98
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_13
timestamp 1626908933
transform 1 0 2688 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_29
timestamp 1626908933
transform 1 0 2688 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_44
timestamp 1626908933
transform 1 0 96 0 -1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_20
timestamp 1626908933
transform 1 0 96 0 -1 6660
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_149
timestamp 1626908933
transform 1 0 3120 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_349
timestamp 1626908933
transform 1 0 3120 0 1 5661
box -32 -32 32 32
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_19
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_79
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_19
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_79
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_12
timestamp 1626908933
transform 1 0 3456 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_73
timestamp 1626908933
transform 1 0 3456 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_30
timestamp 1626908933
transform 1 0 3072 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_14
timestamp 1626908933
transform 1 0 3072 0 -1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_301
timestamp 1626908933
transform 1 0 4080 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_81
timestamp 1626908933
transform 1 0 4080 0 1 5735
box -29 -23 29 23
use M1M2_PR  M1M2_PR_265
timestamp 1626908933
transform 1 0 4272 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_65
timestamp 1626908933
transform 1 0 4272 0 1 5439
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_153
timestamp 1626908933
transform 1 0 3648 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_34
timestamp 1626908933
transform 1 0 3648 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_78
timestamp 1626908933
transform 1 0 3744 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_35
timestamp 1626908933
transform 1 0 3744 0 -1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_302
timestamp 1626908933
transform 1 0 5136 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_300
timestamp 1626908933
transform 1 0 5136 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_82
timestamp 1626908933
transform 1 0 5136 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_80
timestamp 1626908933
transform 1 0 5136 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_230
timestamp 1626908933
transform 1 0 5232 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_30
timestamp 1626908933
transform 1 0 5232 0 1 5661
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_71
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_11
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_71
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_11
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_72
timestamp 1626908933
transform 1 0 4992 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_11
timestamp 1626908933
transform 1 0 4992 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_13
timestamp 1626908933
transform -1 0 4992 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_2
timestamp 1626908933
transform -1 0 4992 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_32
timestamp 1626908933
transform 1 0 5184 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_86
timestamp 1626908933
transform 1 0 5184 0 -1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_260
timestamp 1626908933
transform 1 0 5424 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_258
timestamp 1626908933
transform 1 0 5520 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_40
timestamp 1626908933
transform 1 0 5424 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_38
timestamp 1626908933
transform 1 0 5520 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_228
timestamp 1626908933
transform 1 0 5328 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_28
timestamp 1626908933
transform 1 0 5328 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_120
timestamp 1626908933
transform 1 0 5616 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_320
timestamp 1626908933
transform 1 0 5616 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_13
timestamp 1626908933
transform 1 0 5712 0 1 5513
box -29 -23 29 23
use L1M1_PR  L1M1_PR_233
timestamp 1626908933
transform 1 0 5712 0 1 5513
box -29 -23 29 23
use M1M2_PR  M1M2_PR_10
timestamp 1626908933
transform 1 0 6192 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_210
timestamp 1626908933
transform 1 0 6192 0 1 5587
box -32 -32 32 32
use L1M1_PR  L1M1_PR_10
timestamp 1626908933
transform 1 0 6192 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_230
timestamp 1626908933
transform 1 0 6192 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_142
timestamp 1626908933
transform 1 0 5808 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_362
timestamp 1626908933
transform 1 0 5808 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_18
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_63
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_33
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_152
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_84
timestamp 1626908933
transform 1 0 7536 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_304
timestamp 1626908933
transform 1 0 7536 0 1 5439
box -29 -23 29 23
use M1M2_PR  M1M2_PR_266
timestamp 1626908933
transform 1 0 8112 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_66
timestamp 1626908933
transform 1 0 8112 0 1 5439
box -32 -32 32 32
use L1M1_PR  L1M1_PR_357
timestamp 1626908933
transform 1 0 7728 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_137
timestamp 1626908933
transform 1 0 7728 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_311
timestamp 1626908933
transform 1 0 7920 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_111
timestamp 1626908933
transform 1 0 7920 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_232
timestamp 1626908933
transform 1 0 8112 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_12
timestamp 1626908933
transform 1 0 8112 0 1 5587
box -29 -23 29 23
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_63
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_3
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_63
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_3
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_15
timestamp 1626908933
transform 1 0 7680 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_58
timestamp 1626908933
transform 1 0 7680 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_39
timestamp 1626908933
transform 1 0 5568 0 -1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_15
timestamp 1626908933
transform 1 0 5568 0 -1 6660
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_268
timestamp 1626908933
transform 1 0 8400 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_68
timestamp 1626908933
transform 1 0 8400 0 1 5439
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_71
timestamp 1626908933
transform 1 0 8448 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_10
timestamp 1626908933
transform 1 0 8448 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_63
timestamp 1626908933
transform 1 0 8640 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_9
timestamp 1626908933
transform 1 0 8640 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_48
timestamp 1626908933
transform 1 0 9024 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_5
timestamp 1626908933
transform 1 0 9024 0 -1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_306
timestamp 1626908933
transform 1 0 9264 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_86
timestamp 1626908933
transform 1 0 9264 0 1 5439
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_151
timestamp 1626908933
transform 1 0 9792 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_32
timestamp 1626908933
transform 1 0 9792 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_104
timestamp 1626908933
transform 1 0 9888 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_43
timestamp 1626908933
transform 1 0 9888 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_44
timestamp 1626908933
transform 1 0 0 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_105
timestamp 1626908933
transform 1 0 0 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_99
timestamp 1626908933
transform 1 0 192 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_218
timestamp 1626908933
transform 1 0 192 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_194
timestamp 1626908933
transform 1 0 240 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_394
timestamp 1626908933
transform 1 0 240 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_121
timestamp 1626908933
transform 1 0 144 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_341
timestamp 1626908933
transform 1 0 144 0 1 6327
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_17
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_62
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_93
timestamp 1626908933
transform 1 0 336 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_293
timestamp 1626908933
transform 1 0 336 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_151
timestamp 1626908933
transform 1 0 528 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_371
timestamp 1626908933
transform 1 0 528 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_126
timestamp 1626908933
transform 1 0 720 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_326
timestamp 1626908933
transform 1 0 720 0 1 6401
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_115
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_55
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_115
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_55
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_299
timestamp 1626908933
transform 1 0 1872 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_79
timestamp 1626908933
transform 1 0 1872 0 1 6105
box -29 -23 29 23
use M1M2_PR  M1M2_PR_262
timestamp 1626908933
transform 1 0 1872 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_62
timestamp 1626908933
transform 1 0 1872 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_45
timestamp 1626908933
transform 1 0 2304 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_33
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_21
timestamp 1626908933
transform 1 0 2304 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_9
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_214
timestamp 1626908933
transform 1 0 3312 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_434
timestamp 1626908933
transform 1 0 3312 0 1 6253
box -29 -23 29 23
use M1M2_PR  M1M2_PR_192
timestamp 1626908933
transform 1 0 2928 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_392
timestamp 1626908933
transform 1 0 2928 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_213
timestamp 1626908933
transform 1 0 2928 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_433
timestamp 1626908933
transform 1 0 2928 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_176
timestamp 1626908933
transform 1 0 2832 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_396
timestamp 1626908933
transform 1 0 2832 0 1 6549
box -29 -23 29 23
use M1M2_PR  M1M2_PR_148
timestamp 1626908933
transform 1 0 3120 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_348
timestamp 1626908933
transform 1 0 3120 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_151
timestamp 1626908933
transform 1 0 3312 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_351
timestamp 1626908933
transform 1 0 3312 0 1 6549
box -32 -32 32 32
use L1M1_PR  L1M1_PR_178
timestamp 1626908933
transform 1 0 3216 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_398
timestamp 1626908933
transform 1 0 3216 0 1 6549
box -29 -23 29 23
use M1M2_PR  M1M2_PR_150
timestamp 1626908933
transform 1 0 3312 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_350
timestamp 1626908933
transform 1 0 3312 0 1 6845
box -32 -32 32 32
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_108
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_48
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_108
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_48
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_303
timestamp 1626908933
transform 1 0 4080 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_83
timestamp 1626908933
transform 1 0 4080 0 1 6771
box -29 -23 29 23
use M1M2_PR  M1M2_PR_264
timestamp 1626908933
transform 1 0 4272 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_64
timestamp 1626908933
transform 1 0 4272 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_106
timestamp 1626908933
transform 1 0 4224 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_45
timestamp 1626908933
transform 1 0 4224 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_10
timestamp 1626908933
transform 1 0 4416 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_2
timestamp 1626908933
transform 1 0 4416 0 1 6660
box -38 -49 518 715
use M1M2_PR  M1M2_PR_165
timestamp 1626908933
transform 1 0 4560 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_365
timestamp 1626908933
transform 1 0 4560 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_41
timestamp 1626908933
transform 1 0 4848 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_189
timestamp 1626908933
transform 1 0 4656 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_261
timestamp 1626908933
transform 1 0 4848 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_409
timestamp 1626908933
transform 1 0 4656 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_215
timestamp 1626908933
transform 1 0 4944 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_15
timestamp 1626908933
transform 1 0 4944 0 1 6401
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_219
timestamp 1626908933
transform 1 0 4896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_100
timestamp 1626908933
transform 1 0 4896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_61
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_16
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_231
timestamp 1626908933
transform 1 0 5136 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_31
timestamp 1626908933
transform 1 0 5136 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_150
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_31
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_30
timestamp 1626908933
transform 1 0 5184 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_73
timestamp 1626908933
transform 1 0 5184 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_27
timestamp 1626908933
transform 1 0 5952 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_81
timestamp 1626908933
transform 1 0 5952 0 1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_119
timestamp 1626908933
transform 1 0 5616 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_319
timestamp 1626908933
transform 1 0 5616 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_143
timestamp 1626908933
transform 1 0 5616 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_363
timestamp 1626908933
transform 1 0 5616 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_16
timestamp 1626908933
transform 1 0 6000 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_236
timestamp 1626908933
transform 1 0 6000 0 1 6401
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_41
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_101
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_41
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_101
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use M1M2_PR  M1M2_PR_76
timestamp 1626908933
transform 1 0 7344 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_276
timestamp 1626908933
transform 1 0 7344 0 1 6105
box -32 -32 32 32
use L1M1_PR  L1M1_PR_99
timestamp 1626908933
transform 1 0 7344 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_319
timestamp 1626908933
transform 1 0 7344 0 1 6105
box -29 -23 29 23
use M1M2_PR  M1M2_PR_74
timestamp 1626908933
transform 1 0 7536 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_274
timestamp 1626908933
transform 1 0 7536 0 1 6771
box -32 -32 32 32
use L1M1_PR  L1M1_PR_96
timestamp 1626908933
transform 1 0 7920 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_316
timestamp 1626908933
transform 1 0 7920 0 1 6771
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_30
timestamp 1626908933
transform 1 0 8256 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_149
timestamp 1626908933
transform 1 0 8256 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_27
timestamp 1626908933
transform 1 0 6336 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_3
timestamp 1626908933
transform 1 0 6336 0 1 6660
box -38 -49 1958 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_94
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_34
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_94
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_34
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_57
timestamp 1626908933
transform 1 0 9120 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_3
timestamp 1626908933
transform 1 0 9120 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_53
timestamp 1626908933
transform 1 0 8352 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_10
timestamp 1626908933
transform 1 0 8352 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_29
timestamp 1626908933
transform 1 0 9504 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_101
timestamp 1626908933
transform 1 0 9600 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_148
timestamp 1626908933
transform 1 0 9504 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_220
timestamp 1626908933
transform 1 0 9600 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_15
timestamp 1626908933
transform 1 0 9696 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_60
timestamp 1626908933
transform 1 0 9696 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_46
timestamp 1626908933
transform 1 0 9792 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_107
timestamp 1626908933
transform 1 0 9792 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_102
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_221
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_393
timestamp 1626908933
transform 1 0 48 0 1 7141
box -32 -32 32 32
use M1M2_PR  M1M2_PR_390
timestamp 1626908933
transform 1 0 144 0 1 7511
box -32 -32 32 32
use M1M2_PR  M1M2_PR_193
timestamp 1626908933
transform 1 0 48 0 1 7141
box -32 -32 32 32
use M1M2_PR  M1M2_PR_190
timestamp 1626908933
transform 1 0 144 0 1 7511
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_147
timestamp 1626908933
transform 1 0 0 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_28
timestamp 1626908933
transform 1 0 0 0 -1 7992
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_86
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_26
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_86
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_26
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use L1M1_PR  L1M1_PR_337
timestamp 1626908933
transform 1 0 432 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_117
timestamp 1626908933
transform 1 0 432 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_292
timestamp 1626908933
transform 1 0 336 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_92
timestamp 1626908933
transform 1 0 336 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_107
timestamp 1626908933
transform 1 0 96 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_53
timestamp 1626908933
transform 1 0 96 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_385
timestamp 1626908933
transform 1 0 816 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_165
timestamp 1626908933
transform 1 0 816 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_337
timestamp 1626908933
transform 1 0 912 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_137
timestamp 1626908933
transform 1 0 912 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_432
timestamp 1626908933
transform 1 0 720 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_370
timestamp 1626908933
transform 1 0 624 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_212
timestamp 1626908933
transform 1 0 720 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_150
timestamp 1626908933
transform 1 0 624 0 1 7585
box -29 -23 29 23
use M1M2_PR  M1M2_PR_336
timestamp 1626908933
transform 1 0 912 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_327
timestamp 1626908933
transform 1 0 624 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_136
timestamp 1626908933
transform 1 0 912 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_127
timestamp 1626908933
transform 1 0 624 0 1 7585
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_0
timestamp 1626908933
transform 1 0 480 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_7
timestamp 1626908933
transform 1 0 864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_16
timestamp 1626908933
transform 1 0 480 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_23
timestamp 1626908933
transform 1 0 864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_9
timestamp 1626908933
transform 1 0 1248 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_70
timestamp 1626908933
transform 1 0 1248 0 -1 7992
box -38 -49 230 715
use L1M1_PR  L1M1_PR_164
timestamp 1626908933
transform 1 0 1008 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_384
timestamp 1626908933
transform 1 0 1008 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_309
timestamp 1626908933
transform 1 0 2160 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_89
timestamp 1626908933
transform 1 0 2160 0 1 7215
box -29 -23 29 23
use M1M2_PR  M1M2_PR_271
timestamp 1626908933
transform 1 0 2160 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_270
timestamp 1626908933
transform 1 0 2160 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_71
timestamp 1626908933
transform 1 0 2160 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_70
timestamp 1626908933
transform 1 0 2160 0 1 7437
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_69
timestamp 1626908933
transform 1 0 2208 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_8
timestamp 1626908933
transform 1 0 2208 0 -1 7992
box -38 -49 230 715
use L1M1_PR  L1M1_PR_332
timestamp 1626908933
transform 1 0 2352 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_112
timestamp 1626908933
transform 1 0 2352 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_222
timestamp 1626908933
transform 1 0 2400 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_103
timestamp 1626908933
transform 1 0 2400 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_59
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_14
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_399
timestamp 1626908933
transform 1 0 2736 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_179
timestamp 1626908933
transform 1 0 2736 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_284
timestamp 1626908933
transform 1 0 2640 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_84
timestamp 1626908933
transform 1 0 2640 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_40
timestamp 1626908933
transform 1 0 1440 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_83
timestamp 1626908933
transform 1 0 1440 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_46
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_22
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 1958 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_78
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_18
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_78
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_18
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use M1M2_PR  M1M2_PR_391
timestamp 1626908933
transform 1 0 2928 0 1 7141
box -32 -32 32 32
use M1M2_PR  M1M2_PR_191
timestamp 1626908933
transform 1 0 2928 0 1 7141
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_104
timestamp 1626908933
transform 1 0 4512 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_223
timestamp 1626908933
transform 1 0 4512 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_163
timestamp 1626908933
transform 1 0 4560 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_164
timestamp 1626908933
transform 1 0 4560 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_363
timestamp 1626908933
transform 1 0 4560 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_364
timestamp 1626908933
transform 1 0 4560 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_88
timestamp 1626908933
transform 1 0 4560 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_308
timestamp 1626908933
transform 1 0 4560 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_33
timestamp 1626908933
transform 1 0 4752 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_233
timestamp 1626908933
transform 1 0 4752 0 1 7067
box -32 -32 32 32
use L1M1_PR  L1M1_PR_43
timestamp 1626908933
transform 1 0 4656 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_187
timestamp 1626908933
transform 1 0 4848 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_263
timestamp 1626908933
transform 1 0 4656 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_407
timestamp 1626908933
transform 1 0 4848 0 1 6993
box -29 -23 29 23
use M2M3_PR  M2M3_PR_1
timestamp 1626908933
transform 1 0 4752 0 1 7601
box -33 -37 33 37
use M2M3_PR  M2M3_PR_7
timestamp 1626908933
transform 1 0 4752 0 1 7601
box -33 -37 33 37
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_3
timestamp 1626908933
transform 1 0 4608 0 -1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_15
timestamp 1626908933
transform 1 0 4608 0 -1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_47
timestamp 1626908933
transform 1 0 5280 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_108
timestamp 1626908933
transform 1 0 5280 0 -1 7992
box -38 -49 230 715
use M2M3_PR  M2M3_PR_0
timestamp 1626908933
transform 1 0 5040 0 1 7601
box -33 -37 33 37
use M2M3_PR  M2M3_PR_6
timestamp 1626908933
transform 1 0 5040 0 1 7601
box -33 -37 33 37
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_10
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_70
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_10
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_70
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_105
timestamp 1626908933
transform 1 0 5472 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_224
timestamp 1626908933
transform 1 0 5472 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_15
timestamp 1626908933
transform 1 0 5328 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_235
timestamp 1626908933
transform 1 0 5328 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_318
timestamp 1626908933
transform 1 0 5616 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_118
timestamp 1626908933
transform 1 0 5616 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_80
timestamp 1626908933
transform 1 0 6048 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_26
timestamp 1626908933
transform 1 0 6048 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_1
timestamp 1626908933
transform 1 0 5568 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_12
timestamp 1626908933
transform 1 0 5568 0 -1 7992
box -38 -49 518 715
use M1M2_PR  M1M2_PR_12
timestamp 1626908933
transform 1 0 6480 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_13
timestamp 1626908933
transform 1 0 6480 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_212
timestamp 1626908933
transform 1 0 6480 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_213
timestamp 1626908933
transform 1 0 6480 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_14
timestamp 1626908933
transform 1 0 6768 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_140
timestamp 1626908933
transform 1 0 6384 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_234
timestamp 1626908933
transform 1 0 6768 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_360
timestamp 1626908933
transform 1 0 6384 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_48
timestamp 1626908933
transform 1 0 7200 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_109
timestamp 1626908933
transform 1 0 7200 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_23
timestamp 1626908933
transform 1 0 6432 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_66
timestamp 1626908933
transform 1 0 6432 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_225
timestamp 1626908933
transform 1 0 7392 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_106
timestamp 1626908933
transform 1 0 7392 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_146
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_27
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_58
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_13
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_62
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_2
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_62
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_2
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_14
timestamp 1626908933
transform 1 0 7680 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_57
timestamp 1626908933
transform 1 0 7680 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_68
timestamp 1626908933
transform 1 0 8448 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_7
timestamp 1626908933
transform 1 0 8448 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_62
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_8
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_47
timestamp 1626908933
transform 1 0 9024 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_4
timestamp 1626908933
transform 1 0 9024 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_145
timestamp 1626908933
transform 1 0 9792 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_26
timestamp 1626908933
transform 1 0 9792 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_110
timestamp 1626908933
transform 1 0 9888 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_49
timestamp 1626908933
transform 1 0 9888 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_50
timestamp 1626908933
transform 1 0 0 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_111
timestamp 1626908933
transform 1 0 0 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_107
timestamp 1626908933
transform 1 0 192 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_226
timestamp 1626908933
transform 1 0 192 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_195
timestamp 1626908933
transform 1 0 48 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_395
timestamp 1626908933
transform 1 0 48 0 1 7807
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_12
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_57
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_91
timestamp 1626908933
transform 1 0 336 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_291
timestamp 1626908933
transform 1 0 336 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_116
timestamp 1626908933
transform 1 0 432 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_336
timestamp 1626908933
transform 1 0 432 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_141
timestamp 1626908933
transform 1 0 816 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_341
timestamp 1626908933
transform 1 0 816 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_169
timestamp 1626908933
transform 1 0 816 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_389
timestamp 1626908933
transform 1 0 816 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_215
timestamp 1626908933
transform 1 0 1104 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_435
timestamp 1626908933
transform 1 0 1104 0 1 7733
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_54
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_114
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_54
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_114
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_44
timestamp 1626908933
transform 1 0 2304 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_98
timestamp 1626908933
transform 1 0 2304 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_11
timestamp 1626908933
transform 1 0 2688 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__buf_2  sky130_fd_sc_hs__buf_2_3
timestamp 1626908933
transform 1 0 2688 0 1 7992
box -38 -49 518 715
use M1M2_PR  M1M2_PR_83
timestamp 1626908933
transform 1 0 2640 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_283
timestamp 1626908933
transform 1 0 2640 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_109
timestamp 1626908933
transform 1 0 2640 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_329
timestamp 1626908933
transform 1 0 2640 0 1 7659
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_47
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_23
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_153
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_353
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use L1M1_PR  L1M1_PR_181
timestamp 1626908933
transform 1 0 3024 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_401
timestamp 1626908933
transform 1 0 3024 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_400
timestamp 1626908933
transform 1 0 3312 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_180
timestamp 1626908933
transform 1 0 3312 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_352
timestamp 1626908933
transform 1 0 3312 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_152
timestamp 1626908933
transform 1 0 3312 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_267
timestamp 1626908933
transform 1 0 2928 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_47
timestamp 1626908933
transform 1 0 2928 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_237
timestamp 1626908933
transform 1 0 2928 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_37
timestamp 1626908933
transform 1 0 2928 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_418
timestamp 1626908933
transform 1 0 3120 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_198
timestamp 1626908933
transform 1 0 3120 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_31
timestamp 1626908933
transform 1 0 3168 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_15
timestamp 1626908933
transform 1 0 3168 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_1
timestamp 1626908933
transform 1 0 3552 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_3
timestamp 1626908933
transform 1 0 3552 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_108
timestamp 1626908933
transform 1 0 3936 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_227
timestamp 1626908933
transform 1 0 3936 0 1 7992
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_107
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_47
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_107
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_47
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_311
timestamp 1626908933
transform 1 0 4368 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_91
timestamp 1626908933
transform 1 0 4368 0 1 7881
box -29 -23 29 23
use M1M2_PR  M1M2_PR_372
timestamp 1626908933
transform 1 0 4176 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_172
timestamp 1626908933
transform 1 0 4176 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_269
timestamp 1626908933
transform 1 0 4340 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_49
timestamp 1626908933
transform 1 0 4340 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_2
timestamp 1626908933
transform 1 0 4032 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_14
timestamp 1626908933
transform 1 0 4032 0 1 7992
box -38 -49 710 715
use L1M1_PR  L1M1_PR_310
timestamp 1626908933
transform 1 0 4656 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_90
timestamp 1626908933
transform 1 0 4656 0 1 7881
box -29 -23 29 23
use M1M2_PR  M1M2_PR_235
timestamp 1626908933
transform 1 0 4848 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_234
timestamp 1626908933
transform 1 0 4848 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_35
timestamp 1626908933
transform 1 0 4848 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_34
timestamp 1626908933
transform 1 0 4848 0 1 7807
box -32 -32 32 32
use L1M1_PR  L1M1_PR_266
timestamp 1626908933
transform 1 0 4464 0 1 8335
box -29 -23 29 23
use L1M1_PR  L1M1_PR_237
timestamp 1626908933
transform 1 0 4656 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_46
timestamp 1626908933
transform 1 0 4464 0 1 8335
box -29 -23 29 23
use L1M1_PR  L1M1_PR_17
timestamp 1626908933
transform 1 0 4656 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_239
timestamp 1626908933
transform 1 0 4752 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_39
timestamp 1626908933
transform 1 0 4752 0 1 8177
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_112
timestamp 1626908933
transform 1 0 4704 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_51
timestamp 1626908933
transform 1 0 4704 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_32
timestamp 1626908933
transform 1 0 5040 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_232
timestamp 1626908933
transform 1 0 5040 0 1 7733
box -32 -32 32 32
use L1M1_PR  L1M1_PR_42
timestamp 1626908933
transform 1 0 5040 0 1 7705
box -29 -23 29 23
use L1M1_PR  L1M1_PR_45
timestamp 1626908933
transform 1 0 4902 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_262
timestamp 1626908933
transform 1 0 5040 0 1 7705
box -29 -23 29 23
use L1M1_PR  L1M1_PR_265
timestamp 1626908933
transform 1 0 4902 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_14
timestamp 1626908933
transform 1 0 4944 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_214
timestamp 1626908933
transform 1 0 4944 0 1 8103
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_11
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_56
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_109
timestamp 1626908933
transform 1 0 4896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_228
timestamp 1626908933
transform 1 0 4896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_144
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_25
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_29
timestamp 1626908933
transform 1 0 5184 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_72
timestamp 1626908933
transform 1 0 5184 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_406
timestamp 1626908933
transform 1 0 5616 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_264
timestamp 1626908933
transform 1 0 5712 0 1 7807
box -29 -23 29 23
use L1M1_PR  L1M1_PR_186
timestamp 1626908933
transform 1 0 5616 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_44
timestamp 1626908933
transform 1 0 5712 0 1 7807
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_143
timestamp 1626908933
transform 1 0 5952 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_24
timestamp 1626908933
transform 1 0 5952 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_79
timestamp 1626908933
transform 1 0 6048 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_25
timestamp 1626908933
transform 1 0 6048 0 1 7992
box -38 -49 422 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_100
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_40
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_100
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_40
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_142
timestamp 1626908933
transform 1 0 7200 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_23
timestamp 1626908933
transform 1 0 7200 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_65
timestamp 1626908933
transform 1 0 6432 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_22
timestamp 1626908933
transform 1 0 6432 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_74
timestamp 1626908933
transform 1 0 7296 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_20
timestamp 1626908933
transform 1 0 7296 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_56
timestamp 1626908933
transform 1 0 7680 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_13
timestamp 1626908933
transform 1 0 7680 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_22
timestamp 1626908933
transform 1 0 8448 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_141
timestamp 1626908933
transform 1 0 8448 0 1 7992
box -38 -49 134 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_33
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_93
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_33
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_93
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_3
timestamp 1626908933
transform 1 0 8928 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_46
timestamp 1626908933
transform 1 0 8928 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_7
timestamp 1626908933
transform 1 0 8544 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_61
timestamp 1626908933
transform 1 0 8544 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_229
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_110
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_113
timestamp 1626908933
transform 1 0 9792 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_52
timestamp 1626908933
transform 1 0 9792 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_55
timestamp 1626908933
transform 1 0 9696 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_10
timestamp 1626908933
transform 1 0 9696 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_196
timestamp 1626908933
transform 1 0 48 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_198
timestamp 1626908933
transform 1 0 144 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_396
timestamp 1626908933
transform 1 0 48 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_398
timestamp 1626908933
transform 1 0 144 0 1 9065
box -32 -32 32 32
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_25
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_85
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_25
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_85
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_438
timestamp 1626908933
transform 1 0 1008 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_388
timestamp 1626908933
transform 1 0 912 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_218
timestamp 1626908933
transform 1 0 1008 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_168
timestamp 1626908933
transform 1 0 912 0 1 8917
box -29 -23 29 23
use M1M2_PR  M1M2_PR_340
timestamp 1626908933
transform 1 0 816 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_140
timestamp 1626908933
transform 1 0 816 0 1 8917
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_140
timestamp 1626908933
transform 1 0 1344 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_21
timestamp 1626908933
transform 1 0 1344 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_67
timestamp 1626908933
transform 1 0 1152 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_6
timestamp 1626908933
transform 1 0 1152 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_9
timestamp 1626908933
transform 1 0 768 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_25
timestamp 1626908933
transform 1 0 768 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_42
timestamp 1626908933
transform 1 0 0 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_85
timestamp 1626908933
transform 1 0 0 0 -1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_315
timestamp 1626908933
transform 1 0 2160 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_95
timestamp 1626908933
transform 1 0 2160 0 1 8547
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_139
timestamp 1626908933
transform 1 0 2208 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_20
timestamp 1626908933
transform 1 0 2208 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_114
timestamp 1626908933
transform 1 0 2304 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_53
timestamp 1626908933
transform 1 0 2304 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_54
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_9
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_328
timestamp 1626908933
transform 1 0 2640 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_108
timestamp 1626908933
transform 1 0 2640 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_282
timestamp 1626908933
transform 1 0 2640 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_82
timestamp 1626908933
transform 1 0 2640 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_39
timestamp 1626908933
transform 1 0 1440 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_82
timestamp 1626908933
transform 1 0 1440 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_34
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_10
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_36
timestamp 1626908933
transform 1 0 2928 0 1 8473
box -32 -32 32 32
use M1M2_PR  M1M2_PR_236
timestamp 1626908933
transform 1 0 2928 0 1 8473
box -32 -32 32 32
use L1M1_PR  L1M1_PR_216
timestamp 1626908933
transform 1 0 3408 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_436
timestamp 1626908933
transform 1 0 3408 0 1 8399
box -29 -23 29 23
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_17
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_77
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_17
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_77
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use M1M2_PR  M1M2_PR_145
timestamp 1626908933
transform 1 0 3120 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_345
timestamp 1626908933
transform 1 0 3120 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_173
timestamp 1626908933
transform 1 0 3024 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_393
timestamp 1626908933
transform 1 0 3024 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_93
timestamp 1626908933
transform 1 0 3984 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_94
timestamp 1626908933
transform 1 0 3888 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_313
timestamp 1626908933
transform 1 0 3984 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_314
timestamp 1626908933
transform 1 0 3888 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_73
timestamp 1626908933
transform 1 0 4176 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_273
timestamp 1626908933
transform 1 0 4176 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_72
timestamp 1626908933
transform 1 0 4176 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_272
timestamp 1626908933
transform 1 0 4176 0 1 8769
box -32 -32 32 32
use L1M1_PR  L1M1_PR_92
timestamp 1626908933
transform 1 0 4176 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_312
timestamp 1626908933
transform 1 0 4176 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_362
timestamp 1626908933
transform 1 0 4560 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_162
timestamp 1626908933
transform 1 0 4560 0 1 8991
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_230
timestamp 1626908933
transform 1 0 4512 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_111
timestamp 1626908933
transform 1 0 4512 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_408
timestamp 1626908933
transform 1 0 4656 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_268
timestamp 1626908933
transform 1 0 4752 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_188
timestamp 1626908933
transform 1 0 4656 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_48
timestamp 1626908933
transform 1 0 4752 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_238
timestamp 1626908933
transform 1 0 4752 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_38
timestamp 1626908933
transform 1 0 4752 0 1 8769
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_19
timestamp 1626908933
transform 1 0 5088 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_138
timestamp 1626908933
transform 1 0 5088 0 -1 9324
box -38 -49 134 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_9
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_69
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_9
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_69
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_11
timestamp 1626908933
transform 1 0 4608 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_0
timestamp 1626908933
transform 1 0 4608 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_28
timestamp 1626908933
transform 1 0 5184 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_71
timestamp 1626908933
transform 1 0 5184 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_137
timestamp 1626908933
transform 1 0 5952 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_18
timestamp 1626908933
transform 1 0 5952 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_78
timestamp 1626908933
transform 1 0 6048 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_24
timestamp 1626908933
transform 1 0 6048 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_66
timestamp 1626908933
transform 1 0 7200 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_5
timestamp 1626908933
transform 1 0 7200 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_64
timestamp 1626908933
transform 1 0 6432 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_21
timestamp 1626908933
transform 1 0 6432 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_231
timestamp 1626908933
transform 1 0 7392 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_112
timestamp 1626908933
transform 1 0 7392 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_136
timestamp 1626908933
transform 1 0 7584 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_17
timestamp 1626908933
transform 1 0 7584 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_53
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_8
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_61
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_1
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_61
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_1
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_12
timestamp 1626908933
transform 1 0 7680 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_55
timestamp 1626908933
transform 1 0 7680 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_65
timestamp 1626908933
transform 1 0 8448 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_4
timestamp 1626908933
transform 1 0 8448 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_60
timestamp 1626908933
transform 1 0 8640 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_6
timestamp 1626908933
transform 1 0 8640 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_45
timestamp 1626908933
transform 1 0 9024 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_2
timestamp 1626908933
transform 1 0 9024 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_135
timestamp 1626908933
transform 1 0 9792 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_16
timestamp 1626908933
transform 1 0 9792 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_115
timestamp 1626908933
transform 1 0 9888 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_54
timestamp 1626908933
transform 1 0 9888 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_7
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_52
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_55
timestamp 1626908933
transform 1 0 0 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_116
timestamp 1626908933
transform 1 0 0 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_113
timestamp 1626908933
transform 1 0 192 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_232
timestamp 1626908933
transform 1 0 192 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_197
timestamp 1626908933
transform 1 0 48 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_397
timestamp 1626908933
transform 1 0 48 0 1 9731
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_41
timestamp 1626908933
transform 1 0 768 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_84
timestamp 1626908933
transform 1 0 768 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_52
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_106
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 422 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_113
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_53
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_113
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_53
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_103
timestamp 1626908933
transform 1 0 1536 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_49
timestamp 1626908933
transform 1 0 1536 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_134
timestamp 1626908933
transform 1 0 1920 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_15
timestamp 1626908933
transform 1 0 1920 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_80
timestamp 1626908933
transform 1 0 2016 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_37
timestamp 1626908933
transform 1 0 2016 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_14
timestamp 1626908933
transform 1 0 2784 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_114
timestamp 1626908933
transform 1 0 2880 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_133
timestamp 1626908933
transform 1 0 2784 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_233
timestamp 1626908933
transform 1 0 2880 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_144
timestamp 1626908933
transform 1 0 3120 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_344
timestamp 1626908933
transform 1 0 3120 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_172
timestamp 1626908933
transform 1 0 3120 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_392
timestamp 1626908933
transform 1 0 3120 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_217
timestamp 1626908933
transform 1 0 3216 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_437
timestamp 1626908933
transform 1 0 3216 0 1 9731
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_27
timestamp 1626908933
transform 1 0 2976 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_11
timestamp 1626908933
transform 1 0 2976 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_36
timestamp 1626908933
transform 1 0 3360 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_79
timestamp 1626908933
transform 1 0 3360 0 1 9324
box -38 -49 806 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_106
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_46
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_106
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_46
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_132
timestamp 1626908933
transform 1 0 4128 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_13
timestamp 1626908933
transform 1 0 4128 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_76
timestamp 1626908933
transform 1 0 4224 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_33
timestamp 1626908933
transform 1 0 4224 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_131
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_12
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_70
timestamp 1626908933
transform 1 0 5184 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_27
timestamp 1626908933
transform 1 0 5184 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_51
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_6
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_130
timestamp 1626908933
transform 1 0 5952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_11
timestamp 1626908933
transform 1 0 5952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_77
timestamp 1626908933
transform 1 0 6048 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_23
timestamp 1626908933
transform 1 0 6048 0 1 9324
box -38 -49 422 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_99
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_39
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_99
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_39
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_129
timestamp 1626908933
transform 1 0 7200 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_10
timestamp 1626908933
transform 1 0 7200 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_63
timestamp 1626908933
transform 1 0 6432 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_20
timestamp 1626908933
transform 1 0 6432 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_73
timestamp 1626908933
transform 1 0 7296 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_19
timestamp 1626908933
transform 1 0 7296 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_54
timestamp 1626908933
transform 1 0 7680 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_11
timestamp 1626908933
transform 1 0 7680 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_9
timestamp 1626908933
transform 1 0 8448 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_128
timestamp 1626908933
transform 1 0 8448 0 1 9324
box -38 -49 134 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_32
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_92
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_32
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_92
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1
timestamp 1626908933
transform 1 0 8928 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_44
timestamp 1626908933
transform 1 0 8928 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_5
timestamp 1626908933
transform 1 0 8544 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_59
timestamp 1626908933
transform 1 0 8544 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_234
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_115
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_117
timestamp 1626908933
transform 1 0 9792 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_56
timestamp 1626908933
transform 1 0 9792 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_50
timestamp 1626908933
transform 1 0 9696 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_5
timestamp 1626908933
transform 1 0 9696 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_116
timestamp 1626908933
transform 1 0 192 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_235
timestamp 1626908933
transform 1 0 192 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_176
timestamp 1626908933
transform 1 0 144 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_376
timestamp 1626908933
transform 1 0 144 0 1 10101
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_4
timestamp 1626908933
transform 1 0 288 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_49
timestamp 1626908933
transform 1 0 288 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_8
timestamp 1626908933
transform 1 0 384 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_127
timestamp 1626908933
transform 1 0 384 0 -1 10656
box -38 -49 134 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_24
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_84
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_24
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_84
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_57
timestamp 1626908933
transform 1 0 0 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_118
timestamp 1626908933
transform 1 0 0 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_105
timestamp 1626908933
transform 1 0 480 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_104
timestamp 1626908933
transform 1 0 864 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_51
timestamp 1626908933
transform 1 0 480 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_50
timestamp 1626908933
transform 1 0 864 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_64
timestamp 1626908933
transform 1 0 1248 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_3
timestamp 1626908933
transform 1 0 1248 0 -1 10656
box -38 -49 230 715
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_11
timestamp 1626908933
transform 1 0 1700 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_3
timestamp 1626908933
transform 1 0 1700 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_11
timestamp 1626908933
transform 1 0 1700 0 1 10640
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_3
timestamp 1626908933
transform 1 0 1700 0 1 10640
box -100 -33 100 33
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_126
timestamp 1626908933
transform 1 0 1440 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_7
timestamp 1626908933
transform 1 0 1440 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_102
timestamp 1626908933
transform 1 0 1536 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_48
timestamp 1626908933
transform 1 0 1536 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_119
timestamp 1626908933
transform 1 0 2304 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_58
timestamp 1626908933
transform 1 0 2304 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_101
timestamp 1626908933
transform 1 0 1920 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_47
timestamp 1626908933
transform 1 0 1920 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_96
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_42
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_48
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_76
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_16
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_76
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_16
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_94
timestamp 1626908933
transform 1 0 2976 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_40
timestamp 1626908933
transform 1 0 2976 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_93
timestamp 1626908933
transform 1 0 3360 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_39
timestamp 1626908933
transform 1 0 3360 0 -1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_174
timestamp 1626908933
transform 1 0 3792 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_374
timestamp 1626908933
transform 1 0 3792 0 1 10101
box -32 -32 32 32
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_2
timestamp 1626908933
transform 1 0 4100 0 1 10640
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_10
timestamp 1626908933
transform 1 0 4100 0 1 10640
box -100 -33 100 33
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_2
timestamp 1626908933
transform 1 0 4100 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_10
timestamp 1626908933
transform 1 0 4100 0 1 10633
box -100 -26 100 26
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_38
timestamp 1626908933
transform 1 0 3744 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_92
timestamp 1626908933
transform 1 0 3744 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_2
timestamp 1626908933
transform 1 0 4128 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_63
timestamp 1626908933
transform 1 0 4128 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_125
timestamp 1626908933
transform 1 0 4320 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_6
timestamp 1626908933
transform 1 0 4320 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_91
timestamp 1626908933
transform 1 0 4416 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_37
timestamp 1626908933
transform 1 0 4416 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_236
timestamp 1626908933
transform 1 0 4896 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_124
timestamp 1626908933
transform 1 0 4800 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_117
timestamp 1626908933
transform 1 0 4896 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_5
timestamp 1626908933
transform 1 0 4800 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_47
timestamp 1626908933
transform 1 0 4992 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1626908933
transform 1 0 4992 0 -1 10656
box -38 -49 134 715
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_68
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_8
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_68
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_8
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_123
timestamp 1626908933
transform 1 0 5088 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_4
timestamp 1626908933
transform 1 0 5088 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_85
timestamp 1626908933
transform 1 0 5184 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_31
timestamp 1626908933
transform 1 0 5184 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_122
timestamp 1626908933
transform 1 0 5760 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_3
timestamp 1626908933
transform 1 0 5760 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_62
timestamp 1626908933
transform 1 0 5568 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1
timestamp 1626908933
transform 1 0 5568 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_84
timestamp 1626908933
transform 1 0 5856 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_30
timestamp 1626908933
transform 1 0 5856 0 -1 10656
box -38 -49 422 715
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_9
timestamp 1626908933
transform 1 0 6500 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_1
timestamp 1626908933
transform 1 0 6500 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_9
timestamp 1626908933
transform 1 0 6500 0 1 10640
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_1
timestamp 1626908933
transform 1 0 6500 0 1 10640
box -100 -33 100 33
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_76
timestamp 1626908933
transform 1 0 6240 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_22
timestamp 1626908933
transform 1 0 6240 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_75
timestamp 1626908933
transform 1 0 6624 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_21
timestamp 1626908933
transform 1 0 6624 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_121
timestamp 1626908933
transform 1 0 7008 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_2
timestamp 1626908933
transform 1 0 7008 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_72
timestamp 1626908933
transform 1 0 7104 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_18
timestamp 1626908933
transform 1 0 7104 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_46
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_120
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 134 715
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_0
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA0  hr_16t4_mux_top_VIA0_60
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_0
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use hr_16t4_mux_top_VIA1  hr_16t4_mux_top_VIA1_60
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_15
timestamp 1626908933
transform 1 0 7680 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_69
timestamp 1626908933
transform 1 0 7680 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_68
timestamp 1626908933
transform 1 0 8064 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_14
timestamp 1626908933
transform 1 0 8064 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_119
timestamp 1626908933
transform 1 0 8640 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_0
timestamp 1626908933
transform 1 0 8640 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_61
timestamp 1626908933
transform 1 0 8448 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_0
timestamp 1626908933
transform 1 0 8448 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_58
timestamp 1626908933
transform 1 0 8736 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_4
timestamp 1626908933
transform 1 0 8736 0 -1 10656
box -38 -49 422 715
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_8
timestamp 1626908933
transform 1 0 8900 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA3  hr_16t4_mux_top_VIA3_0
timestamp 1626908933
transform 1 0 8900 0 1 10633
box -100 -26 100 26
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_8
timestamp 1626908933
transform 1 0 8900 0 1 10640
box -100 -33 100 33
use hr_16t4_mux_top_VIA2  hr_16t4_mux_top_VIA2_0
timestamp 1626908933
transform 1 0 8900 0 1 10640
box -100 -33 100 33
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_56
timestamp 1626908933
transform 1 0 9120 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_2
timestamp 1626908933
transform 1 0 9120 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_120
timestamp 1626908933
transform 1 0 9504 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_59
timestamp 1626908933
transform 1 0 9504 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_237
timestamp 1626908933
transform 1 0 9984 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_118
timestamp 1626908933
transform 1 0 9984 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_121
timestamp 1626908933
transform 1 0 9792 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_60
timestamp 1626908933
transform 1 0 9792 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_45
timestamp 1626908933
transform 1 0 9696 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0
timestamp 1626908933
transform 1 0 9696 0 -1 10656
box -38 -49 134 715
<< labels >>
rlabel metal2 s 9922 0 9950 97 4 clk
port 1 nsew
rlabel metal2 s 0 10605 97 10633 4 din[15]
port 2 nsew
rlabel metal2 s 0 9865 97 9893 4 din[14]
port 3 nsew
rlabel metal2 s 0 9125 97 9153 4 din[13]
port 4 nsew
rlabel metal2 s 0 8459 97 8487 4 din[12]
port 5 nsew
rlabel metal2 s 0 7719 97 7747 4 din[11]
port 6 nsew
rlabel metal2 s 0 7053 97 7081 4 din[10]
port 7 nsew
rlabel metal2 s 0 6313 97 6341 4 din[9]
port 8 nsew
rlabel metal2 s 0 5647 97 5675 4 din[8]
port 9 nsew
rlabel metal2 s 0 4907 97 4935 4 din[7]
port 10 nsew
rlabel metal2 s 0 4241 97 4269 4 din[6]
port 11 nsew
rlabel metal2 s 0 3501 97 3529 4 din[5]
port 12 nsew
rlabel metal2 s 0 2835 97 2863 4 din[4]
port 13 nsew
rlabel metal2 s 0 2095 97 2123 4 din[3]
port 14 nsew
rlabel metal2 s 0 1429 97 1457 4 din[2]
port 15 nsew
rlabel metal2 s 0 689 97 717 4 din[1]
port 16 nsew
rlabel metal2 s 0 23 97 51 4 din[0]
port 17 nsew
rlabel metal2 s 130 10559 158 10656 4 rst
port 18 nsew
rlabel metal2 s 130 0 158 97 4 clk_prbs
port 19 nsew
rlabel metal2 s 9983 23 10080 51 4 dout[3]
port 20 nsew
rlabel metal2 s 9983 3575 10080 3603 4 dout[2]
port 21 nsew
rlabel metal2 s 9983 7127 10080 7155 4 dout[1]
port 22 nsew
rlabel metal2 s 9983 10605 10080 10633 4 dout[0]
port 23 nsew
rlabel metal3 s 1600 0 1800 200 4 DVSS:
port 24 nsew
rlabel metal3 s 1600 10456 1800 10656 4 DVSS:
port 24 nsew
rlabel metal3 s 4000 0 4200 200 4 DVSS:
port 24 nsew
rlabel metal3 s 4000 10456 4200 10656 4 DVSS:
port 24 nsew
rlabel metal3 s 6400 0 6600 200 4 DVSS:
port 24 nsew
rlabel metal3 s 6400 10456 6600 10656 4 DVSS:
port 24 nsew
rlabel metal3 s 8800 0 9000 200 4 DVSS:
port 24 nsew
rlabel metal3 s 8800 10456 9000 10656 4 DVSS:
port 24 nsew
rlabel metal1 s 0 -49 98 49 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 -49 10080 49 4 DVSS:
port 24 nsew
rlabel metal1 s 0 1283 98 1381 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 1283 10080 1381 4 DVSS:
port 24 nsew
rlabel metal1 s 0 2615 98 2713 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 2615 10080 2713 4 DVSS:
port 24 nsew
rlabel metal1 s 0 3947 98 4045 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 3947 10080 4045 4 DVSS:
port 24 nsew
rlabel metal1 s 0 5279 98 5377 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 5279 10080 5377 4 DVSS:
port 24 nsew
rlabel metal1 s 0 6611 98 6709 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 6611 10080 6709 4 DVSS:
port 24 nsew
rlabel metal1 s 0 7943 98 8041 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 7943 10080 8041 4 DVSS:
port 24 nsew
rlabel metal1 s 0 9275 98 9373 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 9275 10080 9373 4 DVSS:
port 24 nsew
rlabel metal1 s 0 10607 98 10705 4 DVSS:
port 24 nsew
rlabel metal1 s 9982 10607 10080 10705 4 DVSS:
port 24 nsew
rlabel metal3 s 400 0 600 200 4 DVDD:
port 25 nsew
rlabel metal3 s 400 10456 600 10656 4 DVDD:
port 25 nsew
rlabel metal3 s 2800 0 3000 200 4 DVDD:
port 25 nsew
rlabel metal3 s 2800 10456 3000 10656 4 DVDD:
port 25 nsew
rlabel metal3 s 5200 0 5400 200 4 DVDD:
port 25 nsew
rlabel metal3 s 5200 10456 5400 10656 4 DVDD:
port 25 nsew
rlabel metal3 s 7600 0 7800 200 4 DVDD:
port 25 nsew
rlabel metal3 s 7600 10456 7800 10656 4 DVDD:
port 25 nsew
rlabel metal1 s 0 617 98 715 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 617 10080 715 4 DVDD:
port 25 nsew
rlabel metal1 s 0 1949 98 2047 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 1949 10080 2047 4 DVDD:
port 25 nsew
rlabel metal1 s 0 3281 98 3379 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 3281 10080 3379 4 DVDD:
port 25 nsew
rlabel metal1 s 0 4613 98 4711 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 4613 10080 4711 4 DVDD:
port 25 nsew
rlabel metal1 s 0 5945 98 6043 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 5945 10080 6043 4 DVDD:
port 25 nsew
rlabel metal1 s 0 7277 98 7375 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 7277 10080 7375 4 DVDD:
port 25 nsew
rlabel metal1 s 0 8609 98 8707 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 8609 10080 8707 4 DVDD:
port 25 nsew
rlabel metal1 s 0 9941 98 10039 4 DVDD:
port 25 nsew
rlabel metal1 s 9982 9941 10080 10039 4 DVDD:
port 25 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 26 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 27 nsew
rlabel metal2 s 9936 48 9936 48 4 clk
port 1 nsew
rlabel metal2 s 48 10619 48 10619 4 din[15]
port 2 nsew
rlabel metal2 s 48 9879 48 9879 4 din[14]
port 3 nsew
rlabel metal2 s 48 9139 48 9139 4 din[13]
port 4 nsew
rlabel metal2 s 48 8473 48 8473 4 din[12]
port 5 nsew
rlabel metal2 s 48 7733 48 7733 4 din[11]
port 6 nsew
rlabel metal2 s 48 7067 48 7067 4 din[10]
port 7 nsew
rlabel metal2 s 48 6327 48 6327 4 din[9]
port 8 nsew
rlabel metal2 s 48 5661 48 5661 4 din[8]
port 9 nsew
rlabel metal2 s 48 4921 48 4921 4 din[7]
port 10 nsew
rlabel metal2 s 48 4255 48 4255 4 din[6]
port 11 nsew
rlabel metal2 s 48 3515 48 3515 4 din[5]
port 12 nsew
rlabel metal2 s 48 2849 48 2849 4 din[4]
port 13 nsew
rlabel metal2 s 48 2109 48 2109 4 din[3]
port 14 nsew
rlabel metal2 s 48 1443 48 1443 4 din[2]
port 15 nsew
rlabel metal2 s 48 703 48 703 4 din[1]
port 16 nsew
rlabel metal2 s 48 37 48 37 4 din[0]
port 17 nsew
rlabel metal2 s 144 10607 144 10607 4 rst
port 18 nsew
rlabel metal2 s 144 48 144 48 4 clk_prbs
port 19 nsew
rlabel metal2 s 10031 37 10031 37 4 dout[3]
port 20 nsew
rlabel metal2 s 10031 3589 10031 3589 4 dout[2]
port 21 nsew
rlabel metal2 s 10031 7141 10031 7141 4 dout[1]
port 22 nsew
rlabel metal2 s 10031 10619 10031 10619 4 dout[0]
port 23 nsew
rlabel metal3 s 1700 100 1700 100 4 DVSS:
port 24 nsew
rlabel metal3 s 1700 10556 1700 10556 4 DVSS:
port 24 nsew
rlabel metal3 s 4100 100 4100 100 4 DVSS:
port 24 nsew
rlabel metal3 s 4100 10556 4100 10556 4 DVSS:
port 24 nsew
rlabel metal3 s 6500 100 6500 100 4 DVSS:
port 24 nsew
rlabel metal3 s 6500 10556 6500 10556 4 DVSS:
port 24 nsew
rlabel metal3 s 8900 100 8900 100 4 DVSS:
port 24 nsew
rlabel metal3 s 8900 10556 8900 10556 4 DVSS:
port 24 nsew
rlabel metal1 s 49 0 49 0 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 0 10031 0 4 DVSS:
port 24 nsew
rlabel metal1 s 49 1332 49 1332 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 1332 10031 1332 4 DVSS:
port 24 nsew
rlabel metal1 s 49 2664 49 2664 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 2664 10031 2664 4 DVSS:
port 24 nsew
rlabel metal1 s 49 3996 49 3996 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 3996 10031 3996 4 DVSS:
port 24 nsew
rlabel metal1 s 49 5328 49 5328 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 5328 10031 5328 4 DVSS:
port 24 nsew
rlabel metal1 s 49 6660 49 6660 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 6660 10031 6660 4 DVSS:
port 24 nsew
rlabel metal1 s 49 7992 49 7992 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 7992 10031 7992 4 DVSS:
port 24 nsew
rlabel metal1 s 49 9324 49 9324 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 9324 10031 9324 4 DVSS:
port 24 nsew
rlabel metal1 s 49 10656 49 10656 4 DVSS:
port 24 nsew
rlabel metal1 s 10031 10656 10031 10656 4 DVSS:
port 24 nsew
rlabel metal3 s 500 100 500 100 4 DVDD:
port 25 nsew
rlabel metal3 s 500 10556 500 10556 4 DVDD:
port 25 nsew
rlabel metal3 s 2900 100 2900 100 4 DVDD:
port 25 nsew
rlabel metal3 s 2900 10556 2900 10556 4 DVDD:
port 25 nsew
rlabel metal3 s 5300 100 5300 100 4 DVDD:
port 25 nsew
rlabel metal3 s 5300 10556 5300 10556 4 DVDD:
port 25 nsew
rlabel metal3 s 7700 100 7700 100 4 DVDD:
port 25 nsew
rlabel metal3 s 7700 10556 7700 10556 4 DVDD:
port 25 nsew
rlabel metal1 s 49 666 49 666 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 666 10031 666 4 DVDD:
port 25 nsew
rlabel metal1 s 49 1998 49 1998 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 1998 10031 1998 4 DVDD:
port 25 nsew
rlabel metal1 s 49 3330 49 3330 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 3330 10031 3330 4 DVDD:
port 25 nsew
rlabel metal1 s 49 4662 49 4662 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 4662 10031 4662 4 DVDD:
port 25 nsew
rlabel metal1 s 49 5994 49 5994 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 5994 10031 5994 4 DVDD:
port 25 nsew
rlabel metal1 s 49 7326 49 7326 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 7326 10031 7326 4 DVDD:
port 25 nsew
rlabel metal1 s 49 8658 49 8658 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 8658 10031 8658 4 DVDD:
port 25 nsew
rlabel metal1 s 49 9990 49 9990 4 DVDD:
port 25 nsew
rlabel metal1 s 10031 9990 10031 9990 4 DVDD:
port 25 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 26 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 27 nsew
<< properties >>
string path 126.000 89.725 126.000 119.325 
<< end >>
