magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< locali >>
rect -97 17 96 28
rect -97 -17 -53 17
rect -19 -17 19 17
rect 53 -17 96 17
rect -97 -28 96 -17
<< viali >>
rect -53 -17 -19 17
rect 19 -17 53 17
<< metal1 >>
rect -97 17 96 28
rect -97 -17 -53 17
rect -19 -17 19 17
rect 53 -17 96 17
rect -97 -28 96 -17
<< end >>
