##
## LEF for PtnCells ;
## created by Innovus v19.10-p002_1 on Thu Jun 17 19:36:20 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO digital_top
  CLASS BLOCK ;
  SIZE 550.080000 BY 902.430000 ;
  FOREIGN digital_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 21.1846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.614 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 0.115000 0.485000 0.255000 ;
    END
  END rst
  PIN rst_prbs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.327 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 60.7229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 300.587 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 17.875000 0.485000 18.015000 ;
    END
  END rst_prbs
  PIN inj_error
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.996 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 58.4139 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 289.041 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 36.005000 0.485000 36.145000 ;
    END
  END inj_error
  PIN ref_clk_ext_p
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 154.624 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 235.776 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.155 LAYER met5  ;
    ANTENNAMAXAREACAR 137.714 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 218.253 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 530.080000 572.795000 550.080000 576.795000 ;
    END
  END ref_clk_ext_p
  PIN ref_clk_ext_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.232 LAYER met2  ;
    ANTENNAMAXAREACAR 0.764382 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 0.951165 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0460573 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 530.080000 497.685000 550.080000 501.685000 ;
    END
  END ref_clk_ext_n
  PIN CTL_BUF_N[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0736 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 144.415000 0.485000 144.555000 ;
    END
  END CTL_BUF_N[5]
  PIN CTL_BUF_N[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 2.21991 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.07143 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 126.285000 0.485000 126.425000 ;
    END
  END CTL_BUF_N[4]
  PIN CTL_BUF_N[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 1.37814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 2.72727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 108.155000 0.485000 108.295000 ;
    END
  END CTL_BUF_N[3]
  PIN CTL_BUF_N[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.316 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 52.4017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 258.981 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 90.025000 0.485000 90.165000 ;
    END
  END CTL_BUF_N[2]
  PIN CTL_BUF_N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 1.50087 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 3.34091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 72.265000 0.485000 72.405000 ;
    END
  END CTL_BUF_N[1]
  PIN CTL_BUF_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 1.59329 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 3.80303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 54.135000 0.485000 54.275000 ;
    END
  END CTL_BUF_N[0]
  PIN CTL_BUF_P[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 41.9442 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 206.693 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 252.455000 0.485000 252.595000 ;
    END
  END CTL_BUF_P[5]
  PIN CTL_BUF_P[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.257 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 49.419 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 243.556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 234.325000 0.485000 234.465000 ;
    END
  END CTL_BUF_P[4]
  PIN CTL_BUF_P[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1206 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 58.832 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 291.132 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 216.565000 0.485000 216.705000 ;
    END
  END CTL_BUF_P[3]
  PIN CTL_BUF_P[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 22.324 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.311 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 198.435000 0.485000 198.575000 ;
    END
  END CTL_BUF_P[2]
  PIN CTL_BUF_P[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 33.1229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.587 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 180.305000 0.485000 180.445000 ;
    END
  END CTL_BUF_P[1]
  PIN CTL_BUF_P[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 43.1411 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 212.677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 162.175000 0.485000 162.315000 ;
    END
  END CTL_BUF_P[0]
  PIN osc_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 8.5158 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.947 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 270.585000 0.485000 270.725000 ;
    END
  END osc_en
  PIN aux_osc_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 36.2952 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 177.167 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 288.715000 0.485000 288.855000 ;
    END
  END aux_osc_en
  PIN inj_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 34.1532 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 167.738 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 306.475000 0.485000 306.615000 ;
    END
  END inj_en
  PIN fftl_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 32.7654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 160.799 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 324.605000 0.485000 324.745000 ;
    END
  END fftl_en
  PIN con_perb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.363 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 19.6452 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.9167 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 396.755000 0.485000 396.895000 ;
    END
  END con_perb[3]
  PIN con_perb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0331 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.8561 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 378.625000 0.485000 378.765000 ;
    END
  END con_perb[2]
  PIN con_perb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 32.5411 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 159.677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 360.865000 0.485000 361.005000 ;
    END
  END con_perb[1]
  PIN con_perb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.183 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 33.1654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.799 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 342.735000 0.485000 342.875000 ;
    END
  END con_perb[0]
  PIN div_ratio_half[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.06 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 53.3714 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 263.829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 505.165000 0.485000 505.305000 ;
    END
  END div_ratio_half[5]
  PIN div_ratio_half[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 50.526 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 249.602 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 487.035000 0.485000 487.175000 ;
    END
  END div_ratio_half[4]
  PIN div_ratio_half[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 43.1169 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 212.556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 468.905000 0.485000 469.045000 ;
    END
  END div_ratio_half[3]
  PIN div_ratio_half[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.737 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 36.0805 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 177.374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 451.145000 0.485000 451.285000 ;
    END
  END div_ratio_half[2]
  PIN div_ratio_half[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.586 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 39.129 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.617 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 433.015000 0.485000 433.155000 ;
    END
  END div_ratio_half[1]
  PIN div_ratio_half[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.159 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 42.7836 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.89 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 414.885000 0.485000 415.025000 ;
    END
  END div_ratio_half[0]
  PIN fine_control_avg_window_select[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.982 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 64.5593 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 319.768 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 595.445000 0.485000 595.585000 ;
    END
  END fine_control_avg_window_select[4]
  PIN fine_control_avg_window_select[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.239 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 92.5879 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 458.89 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 577.315000 0.485000 577.455000 ;
    END
  END fine_control_avg_window_select[3]
  PIN fine_control_avg_window_select[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9905 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 48.4351 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.147 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 559.185000 0.485000 559.325000 ;
    END
  END fine_control_avg_window_select[2]
  PIN fine_control_avg_window_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.116 LAYER met2  ;
    ANTENNAMAXAREACAR 8.34476 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.7079 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0460573 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 541.055000 0.485000 541.195000 ;
    END
  END fine_control_avg_window_select[1]
  PIN fine_control_avg_window_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 31.5442 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 154.693 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 523.295000 0.485000 523.435000 ;
    END
  END fine_control_avg_window_select[0]
  PIN fine_con_step_size[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.663 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 87.5022 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 432.95 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 667.595000 0.485000 667.735000 ;
    END
  END fine_con_step_size[3]
  PIN fine_con_step_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.241 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 74.9169 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 371.556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 649.465000 0.485000 649.605000 ;
    END
  END fine_con_step_size[2]
  PIN fine_con_step_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.286 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 60.5957 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 299.95 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 631.335000 0.485000 631.475000 ;
    END
  END fine_con_step_size[1]
  PIN fine_con_step_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.462 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 71.4009 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 353.465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 613.205000 0.485000 613.345000 ;
    END
  END fine_con_step_size[0]
  PIN manual_control_osc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.096 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 49.032 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 242.132 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 902.175000 0.485000 902.315000 ;
    END
  END manual_control_osc[12]
  PIN manual_control_osc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.3265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.246 LAYER met2  ;
    ANTENNAMAXAREACAR 53.8813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 265.435 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.208943 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 884.045000 0.485000 884.185000 ;
    END
  END manual_control_osc[11]
  PIN manual_control_osc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.507 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 29.7169 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 145.556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 865.915000 0.485000 866.055000 ;
    END
  END manual_control_osc[10]
  PIN manual_control_osc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 48.832 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 241.132 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 847.785000 0.485000 847.925000 ;
    END
  END manual_control_osc[9]
  PIN manual_control_osc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.246 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3996 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.5467 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.208943 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 829.655000 0.485000 829.795000 ;
    END
  END manual_control_osc[8]
  PIN manual_control_osc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.563 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 54.2069 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 267.496 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 811.895000 0.485000 812.035000 ;
    END
  END manual_control_osc[7]
  PIN manual_control_osc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.137 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 61.5835 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 304.89 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 793.765000 0.485000 793.905000 ;
    END
  END manual_control_osc[6]
  PIN manual_control_osc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0139 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.9615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 72.7078 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 360.511 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 775.635000 0.485000 775.775000 ;
    END
  END manual_control_osc[5]
  PIN manual_control_osc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4269 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met3  ;
    ANTENNAMAXAREACAR 45.0714 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 225.056 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.395671 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 757.505000 0.485000 757.645000 ;
    END
  END manual_control_osc[4]
  PIN manual_control_osc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.246 LAYER met2  ;
    ANTENNAMAXAREACAR 49.5931 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 243.994 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.208943 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 739.745000 0.485000 739.885000 ;
    END
  END manual_control_osc[3]
  PIN manual_control_osc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 52.1502 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 257.723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 721.615000 0.485000 721.755000 ;
    END
  END manual_control_osc[2]
  PIN manual_control_osc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0226 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.246 LAYER met2  ;
    ANTENNAMAXAREACAR 34.6085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 169.071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.208943 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 703.485000 0.485000 703.625000 ;
    END
  END manual_control_osc[1]
  PIN manual_control_osc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 83.916 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 416.041 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 685.355000 0.485000 685.495000 ;
    END
  END manual_control_osc[0]
  PIN pi1_con[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.728 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 35.2623 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 173.284 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 149.930000 901.945000 150.070000 902.430000 ;
    END
  END pi1_con[3]
  PIN pi1_con[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.7 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 60.9351 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 301.647 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 100.010000 901.945000 100.150000 902.430000 ;
    END
  END pi1_con[2]
  PIN pi1_con[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.92 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 64.6926 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 320.435 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.090000 901.945000 50.230000 902.430000 ;
    END
  END pi1_con[1]
  PIN pi1_con[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.281 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 48.7836 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 240.89 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.650000 901.945000 0.790000 902.430000 ;
    END
  END pi1_con[0]
  PIN pi2_con[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.987 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2937 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.1591 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 349.610000 901.945000 349.750000 902.430000 ;
    END
  END pi2_con[3]
  PIN pi2_con[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.21 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6498 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.0227 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 299.690000 901.945000 299.830000 902.430000 ;
    END
  END pi2_con[2]
  PIN pi2_con[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.21 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0476 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.6477 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 249.770000 901.945000 249.910000 902.430000 ;
    END
  END pi2_con[1]
  PIN pi2_con[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.059 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 51.4199 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 254.071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 199.850000 901.945000 199.990000 902.430000 ;
    END
  END pi2_con[0]
  PIN pi3_con[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.281 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 31.329 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 153.617 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 549.770000 901.945000 549.910000 902.430000 ;
    END
  END pi3_con[3]
  PIN pi3_con[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.37 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.742 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 21.9896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.92 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 499.370000 901.945000 499.510000 902.430000 ;
    END
  END pi3_con[2]
  PIN pi3_con[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 27.1411 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 449.450000 901.945000 449.590000 902.430000 ;
    END
  END pi3_con[1]
  PIN pi3_con[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.987 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5605 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.1705 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 399.530000 901.945000 399.670000 902.430000 ;
    END
  END pi3_con[0]
  PIN pi4_con[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.073 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4787 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.7614 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 147.050000 0.000000 147.190000 0.485000 ;
    END
  END pi4_con[3]
  PIN pi4_con[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.083 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 9.74026 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.6315 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 183.530000 0.000000 183.670000 0.485000 ;
    END
  END pi4_con[2]
  PIN pi4_con[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 7.11266 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.8339 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 220.010000 0.000000 220.150000 0.485000 ;
    END
  END pi4_con[1]
  PIN pi4_con[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.012 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 6.56255 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.2538 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 256.970000 0.000000 257.110000 0.485000 ;
    END
  END pi4_con[0]
  PIN pi5_con[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.763 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 2.95325 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.7381 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.650000 0.000000 0.790000 0.485000 ;
    END
  END pi5_con[3]
  PIN pi5_con[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.663 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 58.2017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 287.981 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 37.130000 0.000000 37.270000 0.485000 ;
    END
  END pi5_con[2]
  PIN pi5_con[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.228 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.231 LAYER met2  ;
    ANTENNAMAXAREACAR 53.3372 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 263.95 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 73.610000 0.000000 73.750000 0.485000 ;
    END
  END pi5_con[1]
  PIN pi5_con[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.404 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.7386 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 110.090000 0.000000 110.230000 0.485000 ;
    END
  END pi5_con[0]
  PIN test_mux_select[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 28.0372 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.023 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 439.850000 0.000000 439.990000 0.485000 ;
    END
  END test_mux_select[3]
  PIN test_mux_select[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.369 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 33.3877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.629 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 476.810000 0.000000 476.950000 0.485000 ;
    END
  END test_mux_select[2]
  PIN test_mux_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.208 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 38.2255 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 184.902 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 513.290000 0.000000 513.430000 0.485000 ;
    END
  END test_mux_select[1]
  PIN test_mux_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.628 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 41.7574 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 204.477 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.111255 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 549.770000 0.000000 549.910000 0.485000 ;
    END
  END test_mux_select[0]
  PIN test_mux_clk_I_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.890000 0.000000 367.030000 0.485000 ;
    END
  END test_mux_clk_I_select[1]
  PIN test_mux_clk_I_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.370000 0.000000 403.510000 0.485000 ;
    END
  END test_mux_clk_I_select[0]
  PIN test_mux_clk_Q_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.450000 0.000000 293.590000 0.485000 ;
    END
  END test_mux_clk_Q_select[1]
  PIN test_mux_clk_Q_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.227 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.924 LAYER met2  ;
    ANTENNAMAXAREACAR 6.99156 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.3674 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0556277 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 330.410000 0.000000 330.550000 0.485000 ;
    END
  END test_mux_clk_Q_select[0]
  PIN dout_p
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 23.1602 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 43.4047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 215.786 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 109.214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 534.365 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.319913 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 415.080000 446.735000 550.080000 452.735000 ;
    END
  END dout_p
  PIN dout_n
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 23.1602 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 36.7687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 182.704 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 LAYER met2  ;
    ANTENNAMAXAREACAR 90.3597 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 440.562 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.222511 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 415.080000 401.965000 550.080000 407.965000 ;
    END
  END dout_n
  PIN test_mux_misc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.6288 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 57.4088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 286.818 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.080000 847.705000 550.080000 851.705000 ;
    END
  END test_mux_misc
  PIN test_mux_clk_Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.221 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.080000 797.755000 550.080000 801.755000 ;
    END
  END test_mux_clk_Q
  PIN test_mux_clk_I
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.994 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.080000 747.805000 550.080000 751.805000 ;
    END
  END test_mux_clk_I
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 400.000000 901.430000 401.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.000000 0.000000 413.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 412.000000 901.430000 413.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.000000 0.000000 425.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.000000 901.430000 425.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.000000 0.000000 437.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 436.000000 901.430000 437.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.000000 0.000000 449.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 448.000000 901.430000 449.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.000000 0.000000 461.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 460.000000 901.430000 461.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.000000 0.000000 473.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 472.000000 901.430000 473.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.000000 0.000000 485.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.000000 901.430000 485.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.000000 0.000000 497.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 496.000000 901.430000 497.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.000000 0.000000 509.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 508.000000 901.430000 509.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.000000 0.000000 521.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 520.000000 901.430000 521.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.000000 0.000000 533.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.000000 901.430000 533.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.000000 0.000000 545.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 544.000000 901.430000 545.000000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 282.240000 900.430000 284.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 262.240000 900.430000 264.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 302.240000 900.430000 304.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 242.240000 900.430000 244.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 322.240000 900.430000 324.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 222.240000 900.430000 224.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 202.240000 900.430000 204.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 182.240000 900.430000 184.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 162.240000 900.430000 164.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 282.240000 0.000000 284.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 262.240000 0.000000 264.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 302.240000 0.000000 304.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 242.240000 0.000000 244.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 322.240000 0.000000 324.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 222.240000 0.000000 224.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 202.240000 0.000000 204.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 182.240000 0.000000 184.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 162.240000 0.000000 164.240000 2.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.240000 901.430000 231.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.160000 901.430000 281.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.160000 901.430000 269.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.160000 901.430000 293.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.160000 901.430000 257.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.160000 901.430000 245.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.080000 901.430000 331.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.080000 901.430000 343.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.240000 901.430000 207.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.080000 901.430000 355.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.240000 901.430000 195.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.080000 901.430000 367.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.240000 901.430000 183.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.080000 901.430000 379.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.240000 901.430000 171.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.240000 901.430000 159.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.160000 0.000000 281.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.160000 0.000000 269.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.160000 0.000000 293.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.160000 0.000000 257.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.160000 0.000000 245.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.080000 0.000000 331.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.080000 0.000000 343.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.240000 0.000000 207.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.080000 0.000000 355.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.240000 0.000000 195.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.080000 0.000000 367.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.240000 0.000000 183.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.080000 0.000000 379.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.240000 0.000000 171.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.240000 0.000000 159.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.320000 901.430000 121.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.320000 901.430000 109.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.320000 901.430000 97.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.320000 901.430000 85.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 901.430000 73.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.320000 0.000000 121.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.320000 0.000000 109.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.320000 0.000000 97.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.320000 0.000000 85.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 0.000000 73.320000 1.000000 ;
    END
  END DVSS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 394.000000 0.000000 395.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.000000 901.430000 395.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.000000 0.000000 407.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 406.000000 901.430000 407.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.000000 0.000000 419.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 418.000000 901.430000 419.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.000000 0.000000 431.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 430.000000 901.430000 431.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.000000 0.000000 443.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 442.000000 901.430000 443.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.000000 0.000000 455.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.000000 901.430000 455.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.000000 0.000000 467.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 466.000000 901.430000 467.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.000000 0.000000 479.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 478.000000 901.430000 479.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.000000 0.000000 491.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 490.000000 901.430000 491.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.000000 0.000000 503.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 502.000000 901.430000 503.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.000000 0.000000 515.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 514.000000 901.430000 515.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.000000 0.000000 527.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 526.000000 901.430000 527.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.000000 0.000000 539.000000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 538.000000 901.430000 539.000000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.240000 901.430000 309.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.240000 901.430000 225.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.160000 901.430000 275.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.160000 901.430000 287.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.160000 901.430000 263.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.160000 901.430000 299.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.160000 901.430000 251.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.160000 901.430000 239.160000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.080000 901.430000 325.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.080000 901.430000 337.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.240000 901.430000 213.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.080000 901.430000 349.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.240000 901.430000 201.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.080000 901.430000 361.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.240000 901.430000 189.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.080000 901.430000 373.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.240000 901.430000 177.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.080000 901.430000 385.080000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.240000 901.430000 165.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.240000 901.430000 153.240000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.160000 0.000000 275.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.160000 0.000000 287.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.160000 0.000000 263.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.160000 0.000000 299.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.160000 0.000000 251.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.160000 0.000000 239.160000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.080000 0.000000 325.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.080000 0.000000 337.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.240000 0.000000 213.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.080000 0.000000 349.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.240000 0.000000 201.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.080000 0.000000 361.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.240000 0.000000 189.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.080000 0.000000 373.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.240000 0.000000 177.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.080000 0.000000 385.080000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.240000 0.000000 165.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.240000 0.000000 153.240000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.320000 901.430000 127.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.320000 901.430000 115.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.320000 901.430000 103.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.320000 901.430000 91.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.320000 901.430000 79.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.320000 901.430000 67.320000 902.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.320000 0.000000 127.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.320000 0.000000 115.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.320000 0.000000 103.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.320000 0.000000 91.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.320000 0.000000 79.320000 1.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.320000 0.000000 67.320000 1.000000 ;
    END
  END DVDD
  PIN AVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 272.240000 900.430000 274.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 292.240000 900.430000 294.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 252.240000 900.430000 254.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 312.240000 900.430000 314.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 232.240000 900.430000 234.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 212.240000 900.430000 214.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 192.240000 900.430000 194.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 172.240000 900.430000 174.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 152.240000 900.430000 154.240000 902.430000 ;
    END
    PORT
      LAYER met5 ;
        RECT 272.240000 0.000000 274.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 292.240000 0.000000 294.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 252.240000 0.000000 254.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 312.240000 0.000000 314.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 232.240000 0.000000 234.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 212.240000 0.000000 214.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 192.240000 0.000000 194.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 172.240000 0.000000 174.240000 2.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 152.240000 0.000000 154.240000 2.000000 ;
    END
  END AVDD
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 550.080000 902.430000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 550.080000 902.430000 ;
    LAYER met2 ;
      RECT 550.050000 901.805000 550.080000 902.430000 ;
      RECT 499.650000 901.805000 549.630000 902.430000 ;
      RECT 449.730000 901.805000 499.230000 902.430000 ;
      RECT 399.810000 901.805000 449.310000 902.430000 ;
      RECT 349.890000 901.805000 399.390000 902.430000 ;
      RECT 299.970000 901.805000 349.470000 902.430000 ;
      RECT 250.050000 901.805000 299.550000 902.430000 ;
      RECT 200.130000 901.805000 249.630000 902.430000 ;
      RECT 150.210000 901.805000 199.710000 902.430000 ;
      RECT 100.290000 901.805000 149.790000 902.430000 ;
      RECT 50.370000 901.805000 99.870000 902.430000 ;
      RECT 0.930000 901.805000 49.950000 902.430000 ;
      RECT 0.000000 901.805000 0.510000 902.035000 ;
      RECT 0.000000 884.325000 550.080000 901.805000 ;
      RECT 0.625000 883.905000 550.080000 884.325000 ;
      RECT 0.000000 866.195000 550.080000 883.905000 ;
      RECT 0.625000 865.775000 550.080000 866.195000 ;
      RECT 0.000000 851.985000 550.080000 865.775000 ;
      RECT 0.000000 848.065000 529.800000 851.985000 ;
      RECT 0.625000 847.645000 529.800000 848.065000 ;
      RECT 0.000000 847.425000 529.800000 847.645000 ;
      RECT 0.000000 829.935000 550.080000 847.425000 ;
      RECT 0.625000 829.515000 550.080000 829.935000 ;
      RECT 0.000000 812.175000 550.080000 829.515000 ;
      RECT 0.625000 811.755000 550.080000 812.175000 ;
      RECT 0.000000 802.035000 550.080000 811.755000 ;
      RECT 0.000000 797.475000 529.800000 802.035000 ;
      RECT 0.000000 794.045000 550.080000 797.475000 ;
      RECT 0.625000 793.625000 550.080000 794.045000 ;
      RECT 0.000000 775.915000 550.080000 793.625000 ;
      RECT 0.625000 775.495000 550.080000 775.915000 ;
      RECT 0.000000 757.785000 550.080000 775.495000 ;
      RECT 0.625000 757.365000 550.080000 757.785000 ;
      RECT 0.000000 752.085000 550.080000 757.365000 ;
      RECT 0.000000 747.525000 529.800000 752.085000 ;
      RECT 0.000000 740.025000 550.080000 747.525000 ;
      RECT 0.625000 739.605000 550.080000 740.025000 ;
      RECT 0.000000 721.895000 550.080000 739.605000 ;
      RECT 0.625000 721.475000 550.080000 721.895000 ;
      RECT 0.000000 703.765000 550.080000 721.475000 ;
      RECT 0.625000 703.345000 550.080000 703.765000 ;
      RECT 0.000000 685.635000 550.080000 703.345000 ;
      RECT 0.625000 685.215000 550.080000 685.635000 ;
      RECT 0.000000 667.875000 550.080000 685.215000 ;
      RECT 0.625000 667.455000 550.080000 667.875000 ;
      RECT 0.000000 649.745000 550.080000 667.455000 ;
      RECT 0.625000 649.325000 550.080000 649.745000 ;
      RECT 0.000000 631.615000 550.080000 649.325000 ;
      RECT 0.625000 631.195000 550.080000 631.615000 ;
      RECT 0.000000 613.485000 550.080000 631.195000 ;
      RECT 0.625000 613.065000 550.080000 613.485000 ;
      RECT 0.000000 595.725000 550.080000 613.065000 ;
      RECT 0.625000 595.305000 550.080000 595.725000 ;
      RECT 0.000000 577.595000 550.080000 595.305000 ;
      RECT 0.625000 577.175000 550.080000 577.595000 ;
      RECT 0.000000 577.075000 550.080000 577.175000 ;
      RECT 0.000000 572.515000 529.800000 577.075000 ;
      RECT 0.000000 559.465000 550.080000 572.515000 ;
      RECT 0.625000 559.045000 550.080000 559.465000 ;
      RECT 0.000000 541.335000 550.080000 559.045000 ;
      RECT 0.625000 540.915000 550.080000 541.335000 ;
      RECT 0.000000 523.575000 550.080000 540.915000 ;
      RECT 0.625000 523.155000 550.080000 523.575000 ;
      RECT 0.000000 505.445000 550.080000 523.155000 ;
      RECT 0.625000 505.025000 550.080000 505.445000 ;
      RECT 0.000000 501.965000 550.080000 505.025000 ;
      RECT 0.000000 497.405000 529.800000 501.965000 ;
      RECT 0.000000 487.315000 550.080000 497.405000 ;
      RECT 0.625000 486.895000 550.080000 487.315000 ;
      RECT 0.000000 469.185000 550.080000 486.895000 ;
      RECT 0.625000 468.765000 550.080000 469.185000 ;
      RECT 0.000000 453.015000 550.080000 468.765000 ;
      RECT 0.000000 451.425000 414.800000 453.015000 ;
      RECT 0.625000 451.005000 414.800000 451.425000 ;
      RECT 0.000000 446.455000 414.800000 451.005000 ;
      RECT 0.000000 433.295000 550.080000 446.455000 ;
      RECT 0.625000 432.875000 550.080000 433.295000 ;
      RECT 0.000000 415.165000 550.080000 432.875000 ;
      RECT 0.625000 414.745000 550.080000 415.165000 ;
      RECT 0.000000 408.245000 550.080000 414.745000 ;
      RECT 0.000000 401.685000 414.800000 408.245000 ;
      RECT 0.000000 397.035000 550.080000 401.685000 ;
      RECT 0.625000 396.615000 550.080000 397.035000 ;
      RECT 0.000000 378.905000 550.080000 396.615000 ;
      RECT 0.625000 378.485000 550.080000 378.905000 ;
      RECT 0.000000 361.145000 550.080000 378.485000 ;
      RECT 0.625000 360.725000 550.080000 361.145000 ;
      RECT 0.000000 343.015000 550.080000 360.725000 ;
      RECT 0.625000 342.595000 550.080000 343.015000 ;
      RECT 0.000000 324.885000 550.080000 342.595000 ;
      RECT 0.625000 324.465000 550.080000 324.885000 ;
      RECT 0.000000 306.755000 550.080000 324.465000 ;
      RECT 0.625000 306.335000 550.080000 306.755000 ;
      RECT 0.000000 288.995000 550.080000 306.335000 ;
      RECT 0.625000 288.575000 550.080000 288.995000 ;
      RECT 0.000000 270.865000 550.080000 288.575000 ;
      RECT 0.625000 270.445000 550.080000 270.865000 ;
      RECT 0.000000 252.735000 550.080000 270.445000 ;
      RECT 0.625000 252.315000 550.080000 252.735000 ;
      RECT 0.000000 234.605000 550.080000 252.315000 ;
      RECT 0.625000 234.185000 550.080000 234.605000 ;
      RECT 0.000000 216.845000 550.080000 234.185000 ;
      RECT 0.625000 216.425000 550.080000 216.845000 ;
      RECT 0.000000 198.715000 550.080000 216.425000 ;
      RECT 0.625000 198.295000 550.080000 198.715000 ;
      RECT 0.000000 180.585000 550.080000 198.295000 ;
      RECT 0.625000 180.165000 550.080000 180.585000 ;
      RECT 0.000000 162.455000 550.080000 180.165000 ;
      RECT 0.625000 162.035000 550.080000 162.455000 ;
      RECT 0.000000 144.695000 550.080000 162.035000 ;
      RECT 0.625000 144.275000 550.080000 144.695000 ;
      RECT 0.000000 126.565000 550.080000 144.275000 ;
      RECT 0.625000 126.145000 550.080000 126.565000 ;
      RECT 0.000000 108.435000 550.080000 126.145000 ;
      RECT 0.625000 108.015000 550.080000 108.435000 ;
      RECT 0.000000 90.305000 550.080000 108.015000 ;
      RECT 0.625000 89.885000 550.080000 90.305000 ;
      RECT 0.000000 72.545000 550.080000 89.885000 ;
      RECT 0.625000 72.125000 550.080000 72.545000 ;
      RECT 0.000000 54.415000 550.080000 72.125000 ;
      RECT 0.625000 53.995000 550.080000 54.415000 ;
      RECT 0.000000 36.285000 550.080000 53.995000 ;
      RECT 0.625000 35.865000 550.080000 36.285000 ;
      RECT 0.000000 18.155000 550.080000 35.865000 ;
      RECT 0.625000 17.735000 550.080000 18.155000 ;
      RECT 0.000000 0.625000 550.080000 17.735000 ;
      RECT 0.000000 0.395000 0.510000 0.625000 ;
      RECT 550.050000 0.000000 550.080000 0.625000 ;
      RECT 513.570000 0.000000 549.630000 0.625000 ;
      RECT 477.090000 0.000000 513.150000 0.625000 ;
      RECT 440.130000 0.000000 476.670000 0.625000 ;
      RECT 403.650000 0.000000 439.710000 0.625000 ;
      RECT 367.170000 0.000000 403.230000 0.625000 ;
      RECT 330.690000 0.000000 366.750000 0.625000 ;
      RECT 293.730000 0.000000 330.270000 0.625000 ;
      RECT 257.250000 0.000000 293.310000 0.625000 ;
      RECT 220.290000 0.000000 256.830000 0.625000 ;
      RECT 183.810000 0.000000 219.870000 0.625000 ;
      RECT 147.330000 0.000000 183.390000 0.625000 ;
      RECT 110.370000 0.000000 146.910000 0.625000 ;
      RECT 73.890000 0.000000 109.950000 0.625000 ;
      RECT 37.410000 0.000000 73.470000 0.625000 ;
      RECT 0.930000 0.000000 36.990000 0.625000 ;
    LAYER met3 ;
      RECT 545.300000 901.130000 550.080000 902.430000 ;
      RECT 539.300000 901.130000 543.700000 902.430000 ;
      RECT 533.300000 901.130000 537.700000 902.430000 ;
      RECT 527.300000 901.130000 531.700000 902.430000 ;
      RECT 521.300000 901.130000 525.700000 902.430000 ;
      RECT 515.300000 901.130000 519.700000 902.430000 ;
      RECT 509.300000 901.130000 513.700000 902.430000 ;
      RECT 503.300000 901.130000 507.700000 902.430000 ;
      RECT 497.300000 901.130000 501.700000 902.430000 ;
      RECT 491.300000 901.130000 495.700000 902.430000 ;
      RECT 485.300000 901.130000 489.700000 902.430000 ;
      RECT 479.300000 901.130000 483.700000 902.430000 ;
      RECT 473.300000 901.130000 477.700000 902.430000 ;
      RECT 467.300000 901.130000 471.700000 902.430000 ;
      RECT 461.300000 901.130000 465.700000 902.430000 ;
      RECT 455.300000 901.130000 459.700000 902.430000 ;
      RECT 449.300000 901.130000 453.700000 902.430000 ;
      RECT 443.300000 901.130000 447.700000 902.430000 ;
      RECT 437.300000 901.130000 441.700000 902.430000 ;
      RECT 431.300000 901.130000 435.700000 902.430000 ;
      RECT 425.300000 901.130000 429.700000 902.430000 ;
      RECT 419.300000 901.130000 423.700000 902.430000 ;
      RECT 413.300000 901.130000 417.700000 902.430000 ;
      RECT 407.300000 901.130000 411.700000 902.430000 ;
      RECT 401.300000 901.130000 405.700000 902.430000 ;
      RECT 395.300000 901.130000 399.700000 902.430000 ;
      RECT 385.380000 901.130000 393.700000 902.430000 ;
      RECT 379.380000 901.130000 383.780000 902.430000 ;
      RECT 373.380000 901.130000 377.780000 902.430000 ;
      RECT 367.380000 901.130000 371.780000 902.430000 ;
      RECT 361.380000 901.130000 365.780000 902.430000 ;
      RECT 355.380000 901.130000 359.780000 902.430000 ;
      RECT 349.380000 901.130000 353.780000 902.430000 ;
      RECT 343.380000 901.130000 347.780000 902.430000 ;
      RECT 337.380000 901.130000 341.780000 902.430000 ;
      RECT 331.380000 901.130000 335.780000 902.430000 ;
      RECT 325.380000 901.130000 329.780000 902.430000 ;
      RECT 309.540000 901.130000 323.780000 902.430000 ;
      RECT 299.460000 901.130000 307.940000 902.430000 ;
      RECT 293.460000 901.130000 297.860000 902.430000 ;
      RECT 287.460000 901.130000 291.860000 902.430000 ;
      RECT 281.460000 901.130000 285.860000 902.430000 ;
      RECT 275.460000 901.130000 279.860000 902.430000 ;
      RECT 269.460000 901.130000 273.860000 902.430000 ;
      RECT 263.460000 901.130000 267.860000 902.430000 ;
      RECT 257.460000 901.130000 261.860000 902.430000 ;
      RECT 251.460000 901.130000 255.860000 902.430000 ;
      RECT 245.460000 901.130000 249.860000 902.430000 ;
      RECT 239.460000 901.130000 243.860000 902.430000 ;
      RECT 231.540000 901.130000 237.860000 902.430000 ;
      RECT 225.540000 901.130000 229.940000 902.430000 ;
      RECT 213.540000 901.130000 223.940000 902.430000 ;
      RECT 207.540000 901.130000 211.940000 902.430000 ;
      RECT 201.540000 901.130000 205.940000 902.430000 ;
      RECT 195.540000 901.130000 199.940000 902.430000 ;
      RECT 189.540000 901.130000 193.940000 902.430000 ;
      RECT 183.540000 901.130000 187.940000 902.430000 ;
      RECT 177.540000 901.130000 181.940000 902.430000 ;
      RECT 171.540000 901.130000 175.940000 902.430000 ;
      RECT 165.540000 901.130000 169.940000 902.430000 ;
      RECT 159.540000 901.130000 163.940000 902.430000 ;
      RECT 153.540000 901.130000 157.940000 902.430000 ;
      RECT 127.620000 901.130000 151.940000 902.430000 ;
      RECT 121.620000 901.130000 126.020000 902.430000 ;
      RECT 115.620000 901.130000 120.020000 902.430000 ;
      RECT 109.620000 901.130000 114.020000 902.430000 ;
      RECT 103.620000 901.130000 108.020000 902.430000 ;
      RECT 97.620000 901.130000 102.020000 902.430000 ;
      RECT 91.620000 901.130000 96.020000 902.430000 ;
      RECT 85.620000 901.130000 90.020000 902.430000 ;
      RECT 79.620000 901.130000 84.020000 902.430000 ;
      RECT 73.620000 901.130000 78.020000 902.430000 ;
      RECT 67.620000 901.130000 72.020000 902.430000 ;
      RECT 0.000000 901.130000 66.020000 902.430000 ;
      RECT 0.000000 1.300000 550.080000 901.130000 ;
      RECT 545.300000 0.000000 550.080000 1.300000 ;
      RECT 539.300000 0.000000 543.700000 1.300000 ;
      RECT 533.300000 0.000000 537.700000 1.300000 ;
      RECT 527.300000 0.000000 531.700000 1.300000 ;
      RECT 521.300000 0.000000 525.700000 1.300000 ;
      RECT 515.300000 0.000000 519.700000 1.300000 ;
      RECT 509.300000 0.000000 513.700000 1.300000 ;
      RECT 503.300000 0.000000 507.700000 1.300000 ;
      RECT 497.300000 0.000000 501.700000 1.300000 ;
      RECT 491.300000 0.000000 495.700000 1.300000 ;
      RECT 485.300000 0.000000 489.700000 1.300000 ;
      RECT 479.300000 0.000000 483.700000 1.300000 ;
      RECT 473.300000 0.000000 477.700000 1.300000 ;
      RECT 467.300000 0.000000 471.700000 1.300000 ;
      RECT 461.300000 0.000000 465.700000 1.300000 ;
      RECT 455.300000 0.000000 459.700000 1.300000 ;
      RECT 449.300000 0.000000 453.700000 1.300000 ;
      RECT 443.300000 0.000000 447.700000 1.300000 ;
      RECT 437.300000 0.000000 441.700000 1.300000 ;
      RECT 431.300000 0.000000 435.700000 1.300000 ;
      RECT 425.300000 0.000000 429.700000 1.300000 ;
      RECT 419.300000 0.000000 423.700000 1.300000 ;
      RECT 413.300000 0.000000 417.700000 1.300000 ;
      RECT 407.300000 0.000000 411.700000 1.300000 ;
      RECT 395.300000 0.000000 405.700000 1.300000 ;
      RECT 385.380000 0.000000 393.700000 1.300000 ;
      RECT 379.380000 0.000000 383.780000 1.300000 ;
      RECT 373.380000 0.000000 377.780000 1.300000 ;
      RECT 367.380000 0.000000 371.780000 1.300000 ;
      RECT 361.380000 0.000000 365.780000 1.300000 ;
      RECT 355.380000 0.000000 359.780000 1.300000 ;
      RECT 349.380000 0.000000 353.780000 1.300000 ;
      RECT 343.380000 0.000000 347.780000 1.300000 ;
      RECT 337.380000 0.000000 341.780000 1.300000 ;
      RECT 331.380000 0.000000 335.780000 1.300000 ;
      RECT 325.380000 0.000000 329.780000 1.300000 ;
      RECT 299.460000 0.000000 323.780000 1.300000 ;
      RECT 293.460000 0.000000 297.860000 1.300000 ;
      RECT 287.460000 0.000000 291.860000 1.300000 ;
      RECT 281.460000 0.000000 285.860000 1.300000 ;
      RECT 275.460000 0.000000 279.860000 1.300000 ;
      RECT 269.460000 0.000000 273.860000 1.300000 ;
      RECT 263.460000 0.000000 267.860000 1.300000 ;
      RECT 257.460000 0.000000 261.860000 1.300000 ;
      RECT 251.460000 0.000000 255.860000 1.300000 ;
      RECT 245.460000 0.000000 249.860000 1.300000 ;
      RECT 239.460000 0.000000 243.860000 1.300000 ;
      RECT 213.540000 0.000000 237.860000 1.300000 ;
      RECT 207.540000 0.000000 211.940000 1.300000 ;
      RECT 201.540000 0.000000 205.940000 1.300000 ;
      RECT 195.540000 0.000000 199.940000 1.300000 ;
      RECT 189.540000 0.000000 193.940000 1.300000 ;
      RECT 183.540000 0.000000 187.940000 1.300000 ;
      RECT 177.540000 0.000000 181.940000 1.300000 ;
      RECT 171.540000 0.000000 175.940000 1.300000 ;
      RECT 165.540000 0.000000 169.940000 1.300000 ;
      RECT 159.540000 0.000000 163.940000 1.300000 ;
      RECT 153.540000 0.000000 157.940000 1.300000 ;
      RECT 127.620000 0.000000 151.940000 1.300000 ;
      RECT 121.620000 0.000000 126.020000 1.300000 ;
      RECT 115.620000 0.000000 120.020000 1.300000 ;
      RECT 109.620000 0.000000 114.020000 1.300000 ;
      RECT 103.620000 0.000000 108.020000 1.300000 ;
      RECT 97.620000 0.000000 102.020000 1.300000 ;
      RECT 91.620000 0.000000 96.020000 1.300000 ;
      RECT 85.620000 0.000000 90.020000 1.300000 ;
      RECT 79.620000 0.000000 84.020000 1.300000 ;
      RECT 73.620000 0.000000 78.020000 1.300000 ;
      RECT 67.620000 0.000000 72.020000 1.300000 ;
      RECT 0.000000 0.000000 66.020000 1.300000 ;
    LAYER met4 ;
      RECT 0.000000 0.000000 550.080000 902.430000 ;
    LAYER met5 ;
      RECT 325.840000 898.830000 550.080000 902.430000 ;
      RECT 315.840000 898.830000 320.640000 902.430000 ;
      RECT 305.840000 898.830000 310.640000 902.430000 ;
      RECT 295.840000 898.830000 300.640000 902.430000 ;
      RECT 285.840000 898.830000 290.640000 902.430000 ;
      RECT 275.840000 898.830000 280.640000 902.430000 ;
      RECT 265.840000 898.830000 270.640000 902.430000 ;
      RECT 255.840000 898.830000 260.640000 902.430000 ;
      RECT 245.840000 898.830000 250.640000 902.430000 ;
      RECT 235.840000 898.830000 240.640000 902.430000 ;
      RECT 225.840000 898.830000 230.640000 902.430000 ;
      RECT 215.840000 898.830000 220.640000 902.430000 ;
      RECT 205.840000 898.830000 210.640000 902.430000 ;
      RECT 195.840000 898.830000 200.640000 902.430000 ;
      RECT 185.840000 898.830000 190.640000 902.430000 ;
      RECT 175.840000 898.830000 180.640000 902.430000 ;
      RECT 165.840000 898.830000 170.640000 902.430000 ;
      RECT 155.840000 898.830000 160.640000 902.430000 ;
      RECT 0.000000 898.830000 150.640000 902.430000 ;
      RECT 0.000000 3.600000 550.080000 898.830000 ;
      RECT 325.840000 0.000000 550.080000 3.600000 ;
      RECT 315.840000 0.000000 320.640000 3.600000 ;
      RECT 305.840000 0.000000 310.640000 3.600000 ;
      RECT 295.840000 0.000000 300.640000 3.600000 ;
      RECT 285.840000 0.000000 290.640000 3.600000 ;
      RECT 275.840000 0.000000 280.640000 3.600000 ;
      RECT 265.840000 0.000000 270.640000 3.600000 ;
      RECT 255.840000 0.000000 260.640000 3.600000 ;
      RECT 245.840000 0.000000 250.640000 3.600000 ;
      RECT 235.840000 0.000000 240.640000 3.600000 ;
      RECT 225.840000 0.000000 230.640000 3.600000 ;
      RECT 215.840000 0.000000 220.640000 3.600000 ;
      RECT 205.840000 0.000000 210.640000 3.600000 ;
      RECT 195.840000 0.000000 200.640000 3.600000 ;
      RECT 185.840000 0.000000 190.640000 3.600000 ;
      RECT 175.840000 0.000000 180.640000 3.600000 ;
      RECT 165.840000 0.000000 170.640000 3.600000 ;
      RECT 155.840000 0.000000 160.640000 3.600000 ;
      RECT 0.000000 0.000000 150.640000 3.600000 ;
  END
END digital_top

END LIBRARY
