magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal2 >>
rect -195 28 195 33
rect -195 -28 -148 28
rect -92 -28 -68 28
rect -12 -28 12 28
rect 68 -28 92 28
rect 148 -28 195 28
rect -195 -33 195 -28
<< via2 >>
rect -148 -28 -92 28
rect -68 -28 -12 28
rect 12 -28 68 28
rect 92 -28 148 28
<< metal3 >>
rect -195 28 195 33
rect -195 -28 -148 28
rect -92 -28 -68 28
rect -12 -28 12 28
rect 68 -28 92 28
rect 148 -28 195 28
rect -195 -33 195 -28
<< end >>
