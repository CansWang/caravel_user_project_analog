magic
tech sky130A
magscale 1 2
timestamp 1624045690
<< error_p >>
rect 1 1 26 610629
rect 511099 587414 511105 587419
rect 511093 587407 511098 587413
rect 511093 587015 511098 587021
rect 511099 587009 511105 587014
rect 510895 567130 510901 567135
rect 510889 567123 510894 567129
rect 510889 566731 510894 566737
rect 510895 566725 510901 566730
use digital_top__user_analog_project_wrapper  digital_top__user_analog_project_wrapper_0
timestamp 1624045690
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
