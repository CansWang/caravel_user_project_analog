magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal3 >>
rect -97 32 96 33
rect -97 -32 -72 32
rect -8 -32 8 32
rect 72 -32 96 32
rect -97 -33 96 -32
<< via3 >>
rect -72 -32 -8 32
rect 8 -32 72 32
<< metal4 >>
rect -97 32 96 33
rect -97 -32 -72 32
rect -8 -32 8 32
rect 72 -32 96 32
rect -97 -33 96 -32
<< end >>
