magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< error_p >>
rect 288 133 289 144
rect 299 99 300 133
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< scpmos >>
rect 84 467 114 551
rect 189 392 289 592
rect 457 368 557 568
rect 628 368 658 592
<< nmoslvt >>
rect 81 74 111 158
rect 253 74 289 158
rect 521 138 557 222
rect 626 74 656 222
<< ndiff >>
rect 405 192 521 222
rect 405 158 413 192
rect 447 158 521 192
rect 28 133 81 158
rect 28 99 36 133
rect 70 99 81 133
rect 28 74 81 99
rect 111 130 253 158
rect 111 96 133 130
rect 167 96 253 130
rect 111 74 253 96
rect 289 133 341 158
rect 405 138 521 158
rect 557 141 626 222
rect 557 138 581 141
rect 289 99 299 133
rect 333 99 341 133
rect 289 74 341 99
rect 573 107 581 138
rect 615 107 626 141
rect 573 74 626 107
rect 656 208 709 222
rect 656 174 667 208
rect 701 174 709 208
rect 656 121 709 174
rect 656 87 667 121
rect 701 87 709 121
rect 656 74 709 87
<< pdiff >>
rect 139 551 189 592
rect 28 529 84 551
rect 28 495 36 529
rect 70 495 84 529
rect 28 467 84 495
rect 114 526 189 551
rect 114 492 131 526
rect 165 492 189 526
rect 114 467 189 492
rect 139 392 189 467
rect 289 529 341 592
rect 573 579 628 592
rect 573 568 581 579
rect 289 495 299 529
rect 333 495 341 529
rect 289 392 341 495
rect 405 422 457 568
rect 405 388 413 422
rect 447 388 457 422
rect 405 368 457 388
rect 557 545 581 568
rect 615 545 628 579
rect 557 471 628 545
rect 557 437 581 471
rect 615 437 628 471
rect 557 368 628 437
rect 658 579 714 592
rect 658 545 672 579
rect 706 545 714 579
rect 658 503 714 545
rect 658 469 672 503
rect 706 469 714 503
rect 658 414 714 469
rect 658 380 672 414
rect 706 380 714 414
rect 658 368 714 380
<< ndiffc >>
rect 413 158 447 192
rect 36 99 70 133
rect 133 96 167 130
rect 299 99 333 133
rect 581 107 615 141
rect 667 174 701 208
rect 667 87 701 121
<< pdiffc >>
rect 36 495 70 529
rect 131 492 165 526
rect 299 495 333 529
rect 413 388 447 422
rect 581 545 615 579
rect 581 437 615 471
rect 672 545 706 579
rect 672 469 706 503
rect 672 380 706 414
<< poly >>
rect 189 592 289 618
rect 84 551 114 577
rect 84 452 114 467
rect 81 304 117 452
rect 457 568 557 594
rect 628 592 658 618
rect 189 344 289 392
rect 189 310 211 344
rect 245 310 289 344
rect 457 326 557 368
rect 628 353 658 368
rect 81 288 147 304
rect 81 254 97 288
rect 131 254 147 288
rect 81 238 147 254
rect 189 276 289 310
rect 189 242 211 276
rect 245 242 289 276
rect 414 310 558 326
rect 625 325 661 353
rect 414 276 430 310
rect 464 276 498 310
rect 532 276 558 310
rect 414 260 558 276
rect 600 309 666 325
rect 600 275 616 309
rect 650 275 666 309
rect 81 158 111 238
rect 189 226 289 242
rect 253 158 289 226
rect 521 222 557 260
rect 600 259 666 275
rect 626 222 656 259
rect 521 112 557 138
rect 81 48 111 74
rect 253 48 289 74
rect 626 48 656 74
<< polycont >>
rect 211 310 245 344
rect 97 254 131 288
rect 211 242 245 276
rect 430 276 464 310
rect 498 276 532 310
rect 616 275 650 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 529 80 545
rect 19 495 36 529
rect 70 495 80 529
rect 19 441 80 495
rect 115 526 181 649
rect 565 579 631 649
rect 565 545 581 579
rect 615 545 631 579
rect 115 492 131 526
rect 165 492 181 526
rect 115 476 181 492
rect 283 529 344 545
rect 283 495 299 529
rect 333 495 344 529
rect 283 479 344 495
rect 19 406 261 441
rect 20 288 146 372
rect 20 254 97 288
rect 131 254 146 288
rect 20 238 146 254
rect 195 344 261 406
rect 195 310 211 344
rect 245 310 261 344
rect 195 276 261 310
rect 195 242 211 276
rect 245 242 261 276
rect 195 204 261 242
rect 19 164 261 204
rect 295 322 344 479
rect 565 471 631 545
rect 397 422 469 438
rect 565 437 581 471
rect 615 437 631 471
rect 565 433 631 437
rect 665 579 748 612
rect 665 545 672 579
rect 706 545 748 579
rect 665 503 748 545
rect 665 469 672 503
rect 706 469 748 503
rect 397 388 413 422
rect 447 399 469 422
rect 665 414 748 469
rect 447 388 631 399
rect 397 365 631 388
rect 582 325 631 365
rect 665 380 672 414
rect 706 380 748 414
rect 665 363 748 380
rect 295 310 548 322
rect 295 276 430 310
rect 464 276 498 310
rect 532 276 548 310
rect 582 309 656 325
rect 19 133 82 164
rect 19 99 36 133
rect 70 99 82 133
rect 295 133 344 276
rect 582 275 616 309
rect 650 275 656 309
rect 582 259 656 275
rect 582 242 631 259
rect 397 208 631 242
rect 690 224 748 363
rect 665 208 748 224
rect 397 192 469 208
rect 397 158 413 192
rect 447 158 469 192
rect 665 174 667 208
rect 701 174 748 208
rect 397 142 469 158
rect 19 61 82 99
rect 117 96 133 130
rect 167 96 183 130
rect 295 127 299 133
rect 117 17 183 96
rect 283 99 299 127
rect 333 99 344 133
rect 283 61 344 99
rect 565 141 631 174
rect 565 107 581 141
rect 615 107 631 141
rect 565 17 631 107
rect 665 121 748 174
rect 665 87 667 121
rect 701 87 748 121
rect 665 71 748 87
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlygate4sd3_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
flabel locali s 703 316 737 350 0 FreeSans 200 0 0 0 X
flabel locali s 703 464 737 498 0 FreeSans 200 0 0 0 X
flabel locali s 703 390 737 424 0 FreeSans 200 0 0 0 X
flabel locali s 703 168 737 202 0 FreeSans 200 0 0 0 X
flabel locali s 703 94 737 128 0 FreeSans 200 0 0 0 X
flabel locali s 703 242 737 276 0 FreeSans 200 0 0 0 X
flabel locali s 703 538 737 572 0 FreeSans 200 0 0 0 X
rlabel comment s 0 0 0 0 4 dlygate4sd3_1
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 384 24 384 24 0 FreeSans 340 0 0 0 VGND
flabel metal1 s 384 641 384 641 0 FreeSans 340 0 0 0 VPWR
flabel locali s 48 259 48 259 0 FreeSans 340 0 0 0 A
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 A
flabel locali s 720 333 720 333 0 FreeSans 200 0 0 0 X
flabel locali s 720 481 720 481 0 FreeSans 200 0 0 0 X
flabel locali s 720 407 720 407 0 FreeSans 200 0 0 0 X
flabel locali s 720 185 720 185 0 FreeSans 200 0 0 0 X
flabel locali s 720 111 720 111 0 FreeSans 200 0 0 0 X
flabel locali s 720 259 720 259 0 FreeSans 200 0 0 0 X
flabel locali s 720 555 720 555 0 FreeSans 200 0 0 0 X
rlabel comment s 0 0 0 0 4 dlygate4sd3_1
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 384 24 384 24 0 FreeSans 340 0 0 0 VGND
flabel metal1 s 384 641 384 641 0 FreeSans 340 0 0 0 VPWR
flabel locali s 48 259 48 259 0 FreeSans 340 0 0 0 A
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 A
flabel locali s 720 333 720 333 0 FreeSans 200 0 0 0 X
flabel locali s 720 481 720 481 0 FreeSans 200 0 0 0 X
flabel locali s 720 407 720 407 0 FreeSans 200 0 0 0 X
flabel locali s 720 185 720 185 0 FreeSans 200 0 0 0 X
flabel locali s 720 111 720 111 0 FreeSans 200 0 0 0 X
flabel locali s 720 259 720 259 0 FreeSans 200 0 0 0 X
flabel locali s 720 555 720 555 0 FreeSans 200 0 0 0 X
<< properties >>
string FIXED_BBOX 0 0 768 666
<< end >>
