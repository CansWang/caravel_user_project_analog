magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal1 >>
rect -83 -26 -58 26
rect -6 -26 6 26
rect 58 -26 83 26
<< via1 >>
rect -58 -26 -6 26
rect 6 -26 58 26
<< metal2 >>
rect -83 -26 -58 26
rect -6 -26 6 26
rect 58 -26 83 26
<< end >>
