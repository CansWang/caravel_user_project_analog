magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 0 0 1248 49
<< scpmos >>
rect 86 368 116 592
rect 280 368 310 592
rect 380 368 410 592
rect 470 368 500 592
rect 765 368 795 592
rect 855 368 885 592
<< nmoslvt >>
rect 82 82 112 230
rect 168 82 198 230
rect 254 82 284 230
rect 340 82 370 230
rect 426 82 456 230
rect 512 82 542 230
rect 598 82 628 230
rect 684 82 714 230
rect 878 82 908 230
rect 964 82 994 230
rect 1050 82 1080 230
rect 1136 82 1166 230
<< ndiff >>
rect 32 164 82 230
rect 27 140 82 164
rect 27 106 37 140
rect 71 106 82 140
rect 27 82 82 106
rect 112 221 168 230
rect 112 187 123 221
rect 157 187 168 221
rect 112 153 168 187
rect 112 119 123 153
rect 157 119 168 153
rect 112 82 168 119
rect 198 140 254 230
rect 198 106 209 140
rect 243 106 254 140
rect 198 82 254 106
rect 284 221 340 230
rect 284 187 295 221
rect 329 187 340 221
rect 284 153 340 187
rect 284 119 295 153
rect 329 119 340 153
rect 284 82 340 119
rect 370 218 426 230
rect 370 184 381 218
rect 415 184 426 218
rect 370 128 426 184
rect 370 94 381 128
rect 415 94 426 128
rect 370 82 426 94
rect 456 221 512 230
rect 456 187 467 221
rect 501 187 512 221
rect 456 153 512 187
rect 456 119 467 153
rect 501 119 512 153
rect 456 82 512 119
rect 542 131 598 230
rect 542 97 553 131
rect 587 97 598 131
rect 542 82 598 97
rect 628 221 684 230
rect 628 187 639 221
rect 673 187 684 221
rect 628 153 684 187
rect 628 119 639 153
rect 673 119 684 153
rect 628 82 684 119
rect 714 164 764 230
rect 714 131 769 164
rect 714 97 725 131
rect 759 97 769 131
rect 714 82 769 97
rect 823 134 878 230
rect 823 100 833 134
rect 867 100 878 134
rect 823 82 878 100
rect 908 218 964 230
rect 908 184 919 218
rect 953 184 964 218
rect 908 128 964 184
rect 908 94 919 128
rect 953 94 964 128
rect 908 82 964 94
rect 994 134 1050 230
rect 994 100 1005 134
rect 1039 100 1050 134
rect 994 82 1050 100
rect 1080 218 1136 230
rect 1080 184 1091 218
rect 1125 184 1136 218
rect 1080 128 1136 184
rect 1080 94 1091 128
rect 1125 94 1136 128
rect 1080 82 1136 94
rect 1166 218 1221 230
rect 1166 184 1177 218
rect 1211 184 1221 218
rect 1166 128 1221 184
rect 1166 94 1177 128
rect 1211 94 1221 128
rect 1166 82 1221 94
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 496 86 546
rect 27 462 39 496
rect 73 462 86 496
rect 27 368 86 462
rect 116 580 280 592
rect 116 546 130 580
rect 164 546 232 580
rect 266 546 280 580
rect 116 510 280 546
rect 116 476 130 510
rect 164 476 232 510
rect 266 476 280 510
rect 116 440 280 476
rect 116 406 130 440
rect 164 406 232 440
rect 266 406 280 440
rect 116 368 280 406
rect 310 580 380 592
rect 310 546 323 580
rect 357 546 380 580
rect 310 508 380 546
rect 310 474 323 508
rect 357 474 380 508
rect 310 368 380 474
rect 410 580 470 592
rect 410 546 423 580
rect 457 546 470 580
rect 410 497 470 546
rect 410 463 423 497
rect 457 463 470 497
rect 410 414 470 463
rect 410 380 423 414
rect 457 380 470 414
rect 410 368 470 380
rect 500 580 765 592
rect 500 546 514 580
rect 548 546 615 580
rect 649 546 717 580
rect 751 546 765 580
rect 500 508 765 546
rect 500 474 514 508
rect 548 474 615 508
rect 649 474 717 508
rect 751 474 765 508
rect 500 368 765 474
rect 795 580 855 592
rect 795 546 808 580
rect 842 546 855 580
rect 795 497 855 546
rect 795 463 808 497
rect 842 463 855 497
rect 795 414 855 463
rect 795 380 808 414
rect 842 380 855 414
rect 795 368 855 380
rect 885 580 1150 592
rect 885 546 899 580
rect 933 546 967 580
rect 1001 546 1035 580
rect 1069 546 1103 580
rect 1137 546 1150 580
rect 885 508 1150 546
rect 885 406 899 508
rect 1137 406 1150 508
rect 885 368 1150 406
<< ndiffc >>
rect 37 106 71 140
rect 123 187 157 221
rect 123 119 157 153
rect 209 106 243 140
rect 295 187 329 221
rect 295 119 329 153
rect 381 184 415 218
rect 381 94 415 128
rect 467 187 501 221
rect 467 119 501 153
rect 553 97 587 131
rect 639 187 673 221
rect 639 119 673 153
rect 725 97 759 131
rect 833 100 867 134
rect 919 184 953 218
rect 919 94 953 128
rect 1005 100 1039 134
rect 1091 184 1125 218
rect 1091 94 1125 128
rect 1177 184 1211 218
rect 1177 94 1211 128
<< pdiffc >>
rect 39 546 73 580
rect 39 462 73 496
rect 130 546 164 580
rect 232 546 266 580
rect 130 476 164 510
rect 232 476 266 510
rect 130 406 164 440
rect 232 406 266 440
rect 323 546 357 580
rect 323 474 357 508
rect 423 546 457 580
rect 423 463 457 497
rect 423 380 457 414
rect 514 546 548 580
rect 615 546 649 580
rect 717 546 751 580
rect 514 474 548 508
rect 615 474 649 508
rect 717 474 751 508
rect 808 546 842 580
rect 808 463 842 497
rect 808 380 842 414
rect 899 546 933 580
rect 967 546 1001 580
rect 1035 546 1069 580
rect 1103 546 1137 580
rect 899 406 1137 508
<< poly >>
rect 86 592 116 618
rect 280 592 310 618
rect 380 592 410 618
rect 470 592 500 618
rect 765 592 795 618
rect 855 592 885 618
rect 86 353 116 368
rect 280 353 310 368
rect 380 353 410 368
rect 470 353 500 368
rect 765 353 795 368
rect 855 353 885 368
rect 83 336 119 353
rect 277 336 313 353
rect 82 320 313 336
rect 377 323 714 353
rect 82 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 313 320
rect 82 275 313 286
rect 426 320 714 323
rect 426 286 442 320
rect 476 286 528 320
rect 562 286 596 320
rect 630 286 664 320
rect 698 286 714 320
rect 82 245 370 275
rect 82 230 112 245
rect 168 230 198 245
rect 254 230 284 245
rect 340 230 370 245
rect 426 270 714 286
rect 426 230 456 270
rect 512 230 542 270
rect 598 230 628 270
rect 684 230 714 270
rect 762 334 798 353
rect 852 334 888 353
rect 762 318 1166 334
rect 762 284 844 318
rect 878 284 912 318
rect 946 284 980 318
rect 1014 284 1048 318
rect 1082 284 1116 318
rect 1150 284 1166 318
rect 762 268 1166 284
rect 878 230 908 268
rect 964 230 994 268
rect 1050 230 1080 268
rect 1136 230 1166 268
rect 82 56 112 82
rect 168 56 198 82
rect 254 56 284 82
rect 340 56 370 82
rect 426 56 456 82
rect 512 56 542 82
rect 598 56 628 82
rect 684 56 714 82
rect 878 56 908 82
rect 964 56 994 82
rect 1050 56 1080 82
rect 1136 56 1166 82
<< polycont >>
rect 121 286 155 320
rect 189 286 223 320
rect 257 286 291 320
rect 442 286 476 320
rect 528 286 562 320
rect 596 286 630 320
rect 664 286 698 320
rect 844 284 878 318
rect 912 284 946 318
rect 980 284 1014 318
rect 1048 284 1082 318
rect 1116 284 1150 318
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 496 89 546
rect 23 462 39 496
rect 73 462 89 496
rect 23 458 89 462
rect 123 580 273 596
rect 123 546 130 580
rect 164 546 232 580
rect 266 546 273 580
rect 123 510 273 546
rect 123 476 130 510
rect 164 476 232 510
rect 266 476 273 510
rect 123 440 273 476
rect 307 580 373 649
rect 307 546 323 580
rect 357 546 373 580
rect 307 508 373 546
rect 307 474 323 508
rect 357 474 373 508
rect 307 458 373 474
rect 407 580 473 596
rect 407 546 423 580
rect 457 546 473 580
rect 407 497 473 546
rect 407 463 423 497
rect 457 463 473 497
rect 123 424 130 440
rect 25 406 130 424
rect 164 406 232 440
rect 266 424 273 440
rect 407 424 473 463
rect 507 580 758 649
rect 507 546 514 580
rect 548 546 615 580
rect 649 546 717 580
rect 751 546 758 580
rect 507 508 758 546
rect 507 474 514 508
rect 548 474 615 508
rect 649 474 717 508
rect 751 474 758 508
rect 507 458 758 474
rect 792 580 858 596
rect 792 546 808 580
rect 842 546 858 580
rect 792 497 858 546
rect 792 463 808 497
rect 842 463 858 497
rect 792 424 858 463
rect 266 414 858 424
rect 266 406 423 414
rect 25 390 423 406
rect 25 236 71 390
rect 407 380 423 390
rect 457 390 808 414
rect 457 380 473 390
rect 407 364 473 380
rect 792 380 808 390
rect 842 380 858 414
rect 892 580 1153 649
rect 892 546 899 580
rect 933 546 967 580
rect 1001 546 1035 580
rect 1069 546 1103 580
rect 1137 546 1153 580
rect 892 508 1153 546
rect 892 406 899 508
rect 1137 406 1153 508
rect 892 390 1153 406
rect 792 364 858 380
rect 105 320 307 356
rect 512 326 743 356
rect 899 326 1223 356
rect 105 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 307 320
rect 105 270 307 286
rect 426 320 743 326
rect 426 286 442 320
rect 476 286 528 320
rect 562 286 596 320
rect 630 286 664 320
rect 698 286 743 320
rect 426 270 743 286
rect 828 318 1223 326
rect 828 284 844 318
rect 878 284 912 318
rect 946 284 980 318
rect 1014 284 1048 318
rect 1082 284 1116 318
rect 1150 284 1223 318
rect 828 268 1223 284
rect 25 221 345 236
rect 25 202 123 221
rect 107 187 123 202
rect 157 202 295 221
rect 157 187 173 202
rect 21 140 71 168
rect 21 106 37 140
rect 107 153 173 187
rect 279 187 295 202
rect 329 187 345 221
rect 107 119 123 153
rect 157 119 173 153
rect 209 140 243 168
rect 21 85 71 106
rect 279 153 345 187
rect 279 119 295 153
rect 329 119 345 153
rect 381 218 415 234
rect 381 128 415 184
rect 209 85 243 106
rect 451 221 1125 234
rect 451 187 467 221
rect 501 187 639 221
rect 673 218 1125 221
rect 673 187 919 218
rect 451 184 919 187
rect 953 184 1091 218
rect 451 153 517 184
rect 451 119 467 153
rect 501 119 517 153
rect 623 153 689 184
rect 551 131 589 150
rect 381 85 415 94
rect 551 97 553 131
rect 587 97 589 131
rect 623 119 639 153
rect 673 119 689 153
rect 723 131 775 150
rect 551 85 589 97
rect 723 97 725 131
rect 759 97 775 131
rect 723 85 775 97
rect 21 51 775 85
rect 817 134 883 150
rect 817 100 833 134
rect 867 100 883 134
rect 817 17 883 100
rect 917 128 955 184
rect 917 94 919 128
rect 953 94 955 128
rect 917 78 955 94
rect 989 134 1055 150
rect 989 100 1005 134
rect 1039 100 1055 134
rect 989 17 1055 100
rect 1091 128 1125 184
rect 1091 78 1125 94
rect 1161 218 1227 234
rect 1161 184 1177 218
rect 1211 184 1227 218
rect 1161 128 1227 184
rect 1161 94 1177 128
rect 1211 94 1227 128
rect 1161 17 1227 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand3_4
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 C
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
rlabel comment s 0 0 0 0 4 nand3_4
flabel pwell s 624 24 624 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 624 641 624 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 624 641 624 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 624 24 624 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 1008 333 1008 333 0 FreeSans 340 0 0 0 C
flabel locali s 1104 333 1104 333 0 FreeSans 340 0 0 0 C
flabel locali s 1200 333 1200 333 0 FreeSans 340 0 0 0 C
flabel locali s 624 333 624 333 0 FreeSans 340 0 0 0 B
flabel locali s 720 333 720 333 0 FreeSans 340 0 0 0 B
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A
flabel locali s 48 259 48 259 0 FreeSans 340 0 0 0 Y
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 Y
rlabel comment s 0 0 0 0 4 nand3_4
flabel pwell s 624 24 624 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 624 641 624 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 624 641 624 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 624 24 624 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 1008 333 1008 333 0 FreeSans 340 0 0 0 C
flabel locali s 1104 333 1104 333 0 FreeSans 340 0 0 0 C
flabel locali s 1200 333 1200 333 0 FreeSans 340 0 0 0 C
flabel locali s 624 333 624 333 0 FreeSans 340 0 0 0 B
flabel locali s 720 333 720 333 0 FreeSans 340 0 0 0 B
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A
flabel locali s 48 259 48 259 0 FreeSans 340 0 0 0 Y
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 1248 666
<< end >>
