magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 0 0 768 49
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 0 617 768 666 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 0 0 768 49 0 FreeSans 200 0 0 0 VGND
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 384 641 384 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 384 641 384 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 384 641 384 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 384 641 384 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 384 641 384 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 384 24 384 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 384 641 384 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_8
flabel metal1 s 384 641 384 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 384 24 384 24 0 FreeSans 200 0 0 0 VGND
<< properties >>
string FIXED_BBOX 0 0 768 666
<< end >>
