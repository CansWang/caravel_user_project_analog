magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 456 368 486 592
rect 546 368 576 592
<< nmoslvt >>
rect 173 80 203 164
rect 344 80 374 164
rect 458 80 488 164
rect 549 80 579 164
<< ndiff >>
rect 27 126 173 164
rect 27 92 39 126
rect 73 92 114 126
rect 148 92 173 126
rect 27 80 173 92
rect 203 141 344 164
rect 203 107 214 141
rect 248 107 299 141
rect 333 107 344 141
rect 203 80 344 107
rect 374 139 458 164
rect 374 105 399 139
rect 433 105 458 139
rect 374 80 458 105
rect 488 139 549 164
rect 488 105 499 139
rect 533 105 549 139
rect 488 80 549 105
rect 579 139 645 164
rect 579 105 599 139
rect 633 105 645 139
rect 579 80 645 105
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 508 86 546
rect 27 474 39 508
rect 73 474 86 508
rect 27 368 86 474
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 504 176 546
rect 116 470 129 504
rect 163 470 176 504
rect 116 424 176 470
rect 116 390 129 424
rect 163 390 176 424
rect 116 368 176 390
rect 206 580 266 592
rect 206 546 219 580
rect 253 546 266 580
rect 206 508 266 546
rect 206 474 219 508
rect 253 474 266 508
rect 206 368 266 474
rect 296 580 356 592
rect 296 546 309 580
rect 343 546 356 580
rect 296 504 356 546
rect 296 470 309 504
rect 343 470 356 504
rect 296 424 356 470
rect 296 390 309 424
rect 343 390 356 424
rect 296 368 356 390
rect 386 580 456 592
rect 386 546 399 580
rect 433 546 456 580
rect 386 508 456 546
rect 386 474 399 508
rect 433 474 456 508
rect 386 368 456 474
rect 486 580 546 592
rect 486 546 499 580
rect 533 546 546 580
rect 486 504 546 546
rect 486 470 499 504
rect 533 470 546 504
rect 486 424 546 470
rect 486 390 499 424
rect 533 390 546 424
rect 486 368 546 390
rect 576 580 645 592
rect 576 546 599 580
rect 633 546 645 580
rect 576 508 645 546
rect 576 474 599 508
rect 633 474 645 508
rect 576 368 645 474
<< ndiffc >>
rect 39 92 73 126
rect 114 92 148 126
rect 214 107 248 141
rect 299 107 333 141
rect 399 105 433 139
rect 499 105 533 139
rect 599 105 633 139
<< pdiffc >>
rect 39 546 73 580
rect 39 474 73 508
rect 129 546 163 580
rect 129 470 163 504
rect 129 390 163 424
rect 219 546 253 580
rect 219 474 253 508
rect 309 546 343 580
rect 309 470 343 504
rect 309 390 343 424
rect 399 546 433 580
rect 399 474 433 508
rect 499 546 533 580
rect 499 470 533 504
rect 499 390 533 424
rect 599 546 633 580
rect 599 474 633 508
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 456 592 486 618
rect 546 592 576 618
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 456 353 486 368
rect 546 353 576 368
rect 83 336 119 353
rect 173 336 209 353
rect 263 336 299 353
rect 353 336 389 353
rect 453 336 489 353
rect 543 336 579 353
rect 83 320 579 336
rect 83 306 189 320
rect 173 286 189 306
rect 223 286 257 320
rect 291 286 325 320
rect 359 286 393 320
rect 427 286 461 320
rect 495 286 579 320
rect 173 270 579 286
rect 173 164 203 270
rect 344 164 374 270
rect 458 164 488 270
rect 549 164 579 270
rect 173 54 203 80
rect 344 54 374 80
rect 458 54 488 80
rect 549 54 579 80
<< polycont >>
rect 189 286 223 320
rect 257 286 291 320
rect 325 286 359 320
rect 393 286 427 320
rect 461 286 495 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 508 73 546
rect 23 474 39 508
rect 23 458 73 474
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 504 179 546
rect 113 470 129 504
rect 163 470 179 504
rect 113 424 179 470
rect 219 580 253 649
rect 219 508 253 546
rect 219 458 253 474
rect 293 580 359 596
rect 293 546 309 580
rect 343 546 359 580
rect 293 504 359 546
rect 293 470 309 504
rect 343 470 359 504
rect 293 424 359 470
rect 399 580 449 649
rect 433 546 449 580
rect 399 508 449 546
rect 433 474 449 508
rect 399 458 449 474
rect 483 580 549 596
rect 483 546 499 580
rect 533 546 549 580
rect 483 504 549 546
rect 483 470 499 504
rect 533 470 549 504
rect 483 424 549 470
rect 583 580 649 649
rect 583 546 599 580
rect 633 546 649 580
rect 583 508 649 546
rect 583 474 599 508
rect 633 474 649 508
rect 583 458 649 474
rect 53 390 129 424
rect 163 390 309 424
rect 343 390 499 424
rect 533 390 647 424
rect 53 236 87 390
rect 121 320 551 356
rect 121 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 286 393 320
rect 427 286 461 320
rect 495 286 551 320
rect 121 270 551 286
rect 601 236 647 390
rect 53 202 647 236
rect 23 126 164 142
rect 23 92 39 126
rect 73 92 114 126
rect 148 92 164 126
rect 23 17 164 92
rect 198 141 349 202
rect 198 107 214 141
rect 248 107 299 141
rect 333 107 349 141
rect 198 91 349 107
rect 383 139 449 168
rect 383 105 399 139
rect 433 105 449 139
rect 383 17 449 105
rect 483 139 549 202
rect 483 105 499 139
rect 533 105 549 139
rect 483 76 549 105
rect 583 139 649 168
rect 583 105 599 139
rect 633 105 649 139
rect 583 17 649 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 clkinv_4
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
rlabel comment s 0 0 0 0 4 clkinv_4
flabel pwell s 336 24 336 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 336 641 336 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 336 641 336 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 336 24 336 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 624 259 624 259 0 FreeSans 340 0 0 0 Y
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A
flabel locali s 336 333 336 333 0 FreeSans 340 0 0 0 A
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 A
flabel locali s 528 333 528 333 0 FreeSans 340 0 0 0 A
rlabel comment s 0 0 0 0 4 clkinv_4
flabel pwell s 336 24 336 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 336 641 336 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 336 641 336 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 336 24 336 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 624 259 624 259 0 FreeSans 340 0 0 0 Y
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A
flabel locali s 336 333 336 333 0 FreeSans 340 0 0 0 A
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 A
flabel locali s 528 333 528 333 0 FreeSans 340 0 0 0 A
rlabel comment s 0 0 0 0 4 clkinv_4
flabel pwell s 336 24 336 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 336 641 336 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 336 641 336 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 336 24 336 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 624 259 624 259 0 FreeSans 340 0 0 0 Y
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A
flabel locali s 336 333 336 333 0 FreeSans 340 0 0 0 A
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 A
flabel locali s 528 333 528 333 0 FreeSans 340 0 0 0 A
rlabel comment s 0 0 0 0 4 clkinv_4
flabel pwell s 336 24 336 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 336 641 336 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 336 641 336 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 336 24 336 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 624 259 624 259 0 FreeSans 340 0 0 0 Y
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A
flabel locali s 336 333 336 333 0 FreeSans 340 0 0 0 A
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 A
flabel locali s 528 333 528 333 0 FreeSans 340 0 0 0 A
<< properties >>
string FIXED_BBOX 0 0 672 666
<< end >>
