magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal1 >>
rect -292 26 292 49
rect -292 -26 -282 26
rect -230 -26 -218 26
rect -166 -26 -154 26
rect -102 -26 -90 26
rect -38 -26 -26 26
rect 26 -26 38 26
rect 90 -26 102 26
rect 154 -26 166 26
rect 218 -26 230 26
rect 282 -26 292 26
rect -292 -49 292 -26
<< via1 >>
rect -282 -26 -230 26
rect -218 -26 -166 26
rect -154 -26 -102 26
rect -90 -26 -38 26
rect -26 -26 26 26
rect 38 -26 90 26
rect 102 -26 154 26
rect 166 -26 218 26
rect 230 -26 282 26
<< metal2 >>
rect -292 26 292 49
rect -292 -26 -282 26
rect -230 -26 -218 26
rect -166 -26 -154 26
rect -102 -26 -90 26
rect -38 -26 -26 26
rect 26 -26 38 26
rect 90 -26 102 26
rect 154 -26 166 26
rect 218 -26 230 26
rect 282 -26 292 26
rect -292 -49 292 -26
<< end >>
