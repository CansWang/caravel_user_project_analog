magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< error_s >>
rect 1118 13431 1119 13476
rect 2270 13431 2271 13476
rect 3518 13431 3519 13476
rect 4574 13431 4575 13476
rect 5438 13431 5439 13476
rect 7166 13431 7167 13476
rect 8414 13431 8415 13476
rect 9566 13431 9567 13476
rect 10814 13431 10815 13476
rect 12062 13431 12063 13476
rect 13214 13431 13215 13476
rect 446 13175 447 13220
rect 1694 13175 1695 13220
rect 2942 13175 2943 13220
rect 4094 13175 4095 13220
rect 5918 13175 5919 13220
rect 7070 13175 7071 13220
rect 10814 13175 10815 13220
rect 12062 13175 12063 13220
rect 13310 13175 13311 13220
rect 1118 12099 1119 12144
rect 2270 12099 2271 12144
rect 3134 12099 3135 12144
rect 7742 12099 7743 12144
rect 8990 12099 8991 12144
rect 10814 12099 10815 12144
rect 12062 12099 12063 12144
rect 13214 12099 13215 12144
rect 446 11843 447 11888
rect 1694 11843 1695 11888
rect 2942 11843 2943 11888
rect 4094 11843 4095 11888
rect 5918 11843 5919 11888
rect 10814 11843 10815 11888
rect 12062 11843 12063 11888
rect 13310 11843 13311 11888
rect 1118 10767 1119 10812
rect 1886 10767 1887 10812
rect 4574 10767 4575 10812
rect 10814 10767 10815 10812
rect 12062 10767 12063 10812
rect 13214 10767 13215 10812
rect 446 10511 447 10556
rect 5918 10511 5919 10556
rect 7070 10511 7071 10556
rect 830 9435 831 9480
rect 5726 9435 5727 9480
rect 446 9179 447 9224
rect 1694 9179 1695 9224
rect 9374 9179 9375 9224
rect 12062 9179 12063 9224
rect 926 8103 927 8148
rect 3518 8103 3519 8148
rect 4574 8103 4575 8148
rect 5534 8103 5535 8148
rect 446 7847 447 7892
rect 2942 7847 2943 7892
rect 5918 7847 5919 7892
rect 7070 7847 7071 7892
rect 8222 7847 8223 7892
rect 10142 7847 10143 7892
rect 12926 7847 12927 7892
rect 734 6771 735 6816
rect 3518 6771 3519 6816
rect 5438 6771 5439 6816
rect 446 6515 447 6560
rect 5054 6515 5055 6560
rect 8414 6515 8415 6560
rect 9662 6515 9663 6560
rect 12062 6515 12063 6560
rect 13214 6515 13215 6560
rect 1118 5439 1119 5484
rect 10814 5439 10815 5484
rect 350 5183 351 5228
rect 2078 5183 2079 5228
rect 10718 4107 10719 4152
rect 446 3851 447 3896
rect 2078 3851 2079 3896
rect 4862 3851 4863 3896
rect 7070 3851 7071 3896
rect 11486 3851 11487 3896
rect 1118 2775 1119 2820
rect 7742 2775 7743 2820
rect 8990 2775 8991 2820
rect 446 2519 447 2564
rect 1694 2519 1695 2564
rect 2942 2519 2943 2564
rect 3902 2519 3903 2564
rect 13310 2519 13311 2564
rect 1118 1443 1119 1488
rect 5438 1443 5439 1488
rect 446 1187 447 1232
rect 1694 1187 1695 1232
rect 2942 1187 2943 1232
rect 3710 1187 3711 1232
rect 6590 1187 6591 1232
rect 13310 1187 13311 1232
rect 1118 111 1119 156
rect 2078 111 2079 156
rect 7934 111 7935 156
rect 9566 111 9567 156
rect 12062 111 12063 156
rect 13310 111 13311 156
<< locali >>
rect 9264 13044 9377 13078
rect 9343 12970 9377 13044
rect 5119 12338 5153 12412
rect 3487 12264 3521 12338
rect 4752 12304 5153 12338
rect 5695 12264 5729 12560
rect 6576 12304 6689 12338
rect 3487 12230 3600 12264
rect 5616 12230 5729 12264
rect 4447 11860 4656 11894
rect 8575 11860 8688 11894
rect 4447 11712 4481 11860
rect 10015 11746 10049 11894
rect 4543 11672 4577 11746
rect 9936 11712 10049 11746
rect 4543 11638 4656 11672
rect 3103 10414 3137 10562
rect 12415 10414 12449 10562
rect 3024 10380 3137 10414
rect 12336 10380 12449 10414
rect 2623 9600 2657 9896
rect 10495 9600 10529 9748
rect 2544 9566 2657 9600
rect 10416 9566 10529 9600
rect 8095 9082 8129 9156
rect 6079 9048 6288 9082
rect 7711 9048 7824 9082
rect 8016 9048 8129 9082
rect 6079 8900 6113 9048
rect 7711 8752 7745 9048
rect 6655 8308 6768 8342
rect 8287 8308 8400 8342
rect 10399 8268 10433 8416
rect 11071 8342 11105 8564
rect 11071 8308 11184 8342
rect 10320 8234 10433 8268
rect 1279 7864 1392 7898
rect 1279 7420 1313 7864
rect 9727 7750 9761 7898
rect 8880 7716 8993 7750
rect 9648 7716 9761 7750
rect 8959 7568 8993 7716
rect 4447 6936 4481 7158
rect 7423 6976 7536 7010
rect 4368 6902 4481 6936
rect 5791 6902 5904 6936
rect 8959 6902 9072 6936
rect 8959 6828 8993 6902
rect 1471 6532 1584 6566
rect 895 6384 1008 6418
rect 895 6162 929 6384
rect 1471 6088 1505 6532
rect 2160 6458 2273 6492
rect 13567 6384 13680 6418
rect 13567 6088 13601 6384
rect 4752 5570 4865 5604
rect 4831 5496 4865 5570
rect 6079 5570 6192 5604
rect 6079 5422 6113 5570
rect 10399 5012 10433 5234
rect 10320 4978 10433 5012
rect 2719 4346 2753 4494
rect 2640 4312 2753 4346
rect 5599 3754 5633 3902
rect 5520 3720 5633 3754
rect 6175 3720 6288 3754
rect 6480 3720 6593 3754
rect 6175 3424 6209 3720
rect 6559 3424 6593 3720
rect 10207 3680 10241 3828
rect 10128 3646 10241 3680
rect 13488 1574 13601 1608
rect 13567 1500 13601 1574
rect 8959 982 9264 1016
rect 7135 128 7169 498
rect 9055 350 9089 572
rect 8976 316 9089 350
rect 10687 276 10721 572
rect 10687 242 10800 276
rect 7056 94 7169 128
<< metal1 >>
rect 0 14603 14016 14701
rect 4834 14379 6014 14407
rect 6178 14379 8606 14407
rect 418 14231 4670 14259
rect 418 14185 446 14231
rect 226 14157 446 14185
rect 4642 14185 4670 14231
rect 4642 14157 8414 14185
rect 6009 14083 6096 14111
rect 0 13937 14016 14035
rect 5410 13713 6206 13741
rect 6082 13639 6206 13667
rect 6082 13417 6494 13445
rect 0 13271 14016 13369
rect 5218 13195 5438 13223
rect 9250 13121 11678 13149
rect 4953 13047 5040 13075
rect 5145 13047 5232 13075
rect 8985 13047 9072 13075
rect 9250 13001 9278 13121
rect 226 12973 4862 13001
rect 4834 12927 4862 12973
rect 5314 12973 6878 13001
rect 7906 12973 8414 13001
rect 8505 12973 8592 13001
rect 8674 12973 9278 13001
rect 9346 12973 9566 13001
rect 5314 12927 5342 12973
rect 8386 12927 8414 12973
rect 9538 12927 9566 12973
rect 11746 12973 12734 13001
rect 11746 12927 11774 12973
rect 4834 12899 5342 12927
rect 7906 12899 8222 12927
rect 8386 12899 8510 12927
rect 9538 12899 11774 12927
rect 8194 12853 8222 12899
rect 8194 12825 9182 12853
rect 7522 12751 7838 12779
rect 0 12605 14016 12703
rect 5698 12529 5918 12557
rect 5890 12520 5918 12529
rect 9346 12529 9566 12557
rect 10882 12529 11102 12557
rect 5890 12492 6494 12520
rect 6466 12483 6494 12492
rect 6466 12455 7742 12483
rect 7714 12409 7742 12455
rect 9346 12409 9374 12529
rect 3682 12381 4478 12409
rect 5122 12381 6302 12409
rect 7714 12381 9374 12409
rect 11074 12409 11102 12529
rect 12514 12529 12734 12557
rect 12514 12409 12542 12529
rect 11074 12381 12542 12409
rect 898 12307 3518 12335
rect 4450 12307 5534 12335
rect 6082 12307 6302 12335
rect 6658 12307 6974 12335
rect 7042 12307 7550 12335
rect 3778 12233 3902 12261
rect 5337 12233 5424 12261
rect 7906 12159 8414 12187
rect 7906 12113 7934 12159
rect 7042 12085 7358 12113
rect 7714 12085 7934 12113
rect 8386 12113 8414 12159
rect 8386 12085 8606 12113
rect 0 11939 14016 12037
rect 226 11863 638 11891
rect 610 11817 638 11863
rect 6178 11863 6398 11891
rect 6850 11863 7646 11891
rect 8386 11863 8606 11891
rect 10018 11863 10718 11891
rect 6178 11854 6206 11863
rect 1474 11826 6206 11854
rect 1474 11817 1502 11826
rect 610 11789 1502 11817
rect 226 11715 446 11743
rect 418 11595 446 11715
rect 4258 11715 4478 11743
rect 4546 11715 5438 11743
rect 5602 11715 9086 11743
rect 9250 11715 9758 11743
rect 4258 11669 4286 11715
rect 5602 11669 5630 11715
rect 1666 11641 4286 11669
rect 1666 11595 1694 11641
rect 418 11567 1694 11595
rect 4930 11521 4958 11669
rect 5026 11641 5630 11669
rect 6466 11641 6590 11669
rect 6658 11595 6686 11669
rect 6754 11641 6782 11715
rect 7641 11641 7728 11669
rect 7810 11641 7934 11669
rect 8002 11641 8030 11715
rect 8697 11641 8784 11669
rect 8866 11641 8990 11669
rect 9058 11641 9086 11715
rect 7810 11595 7838 11641
rect 8866 11595 8894 11641
rect 6658 11567 11102 11595
rect 5122 11530 5918 11558
rect 5122 11521 5150 11530
rect 1858 11493 5150 11521
rect 5890 11521 5918 11530
rect 6658 11521 6686 11567
rect 5890 11493 6686 11521
rect 7138 11456 7838 11484
rect 7138 11447 7166 11456
rect 5218 11419 5822 11447
rect 6946 11419 7166 11447
rect 7810 11447 7838 11456
rect 7810 11419 8030 11447
rect 8121 11419 8208 11447
rect 9250 11419 9470 11447
rect 9634 11419 9854 11447
rect 0 11273 14016 11371
rect 2818 11197 3614 11225
rect 3586 11188 3614 11197
rect 4930 11197 5150 11225
rect 6562 11197 7166 11225
rect 8770 11197 9182 11225
rect 4930 11188 4958 11197
rect 3586 11160 4958 11188
rect 7138 11188 7166 11197
rect 7138 11160 7838 11188
rect 7810 11151 7838 11160
rect 7810 11123 8414 11151
rect 8386 11077 8414 11123
rect 9058 11123 9278 11151
rect 9058 11077 9086 11123
rect 8386 11049 9086 11077
rect 2530 10975 3422 11003
rect 3586 10975 7646 11003
rect 8002 10975 8222 11003
rect 2530 10929 2558 10975
rect 1474 10901 2174 10929
rect 2338 10901 2558 10929
rect 3394 10929 3422 10975
rect 3394 10901 3806 10929
rect 5721 10901 5808 10929
rect 10882 10901 12542 10929
rect 1474 10781 1502 10901
rect 1282 10753 1502 10781
rect 2146 10781 2174 10901
rect 10882 10855 10910 10901
rect 10690 10827 10910 10855
rect 12514 10855 12542 10901
rect 12514 10827 12734 10855
rect 2626 10790 4670 10818
rect 2626 10781 2654 10790
rect 2146 10753 2654 10781
rect 4642 10781 4670 10790
rect 4642 10753 4862 10781
rect 0 10607 14016 10705
rect 226 10531 446 10559
rect 418 10485 446 10531
rect 994 10531 1214 10559
rect 1762 10531 1982 10559
rect 3106 10531 3230 10559
rect 5314 10531 5534 10559
rect 8578 10531 9182 10559
rect 12418 10531 12638 10559
rect 994 10485 1022 10531
rect 1954 10522 1982 10531
rect 12610 10522 12638 10531
rect 13282 10531 13502 10559
rect 13282 10522 13310 10531
rect 1954 10494 2846 10522
rect 12610 10494 13310 10522
rect 418 10457 1022 10485
rect 2818 10485 2846 10494
rect 2818 10457 2942 10485
rect 2914 10411 2942 10457
rect 11362 10411 11390 10485
rect 1666 10383 2846 10411
rect 2914 10383 3998 10411
rect 7929 10383 8016 10411
rect 9442 10383 10046 10411
rect 11362 10383 12350 10411
rect 12898 10383 13022 10411
rect 13186 10383 13310 10411
rect 1209 10309 1296 10337
rect 1474 10189 1502 10337
rect 1570 10309 1886 10337
rect 3513 10309 3600 10337
rect 7545 10309 9662 10337
rect 1858 10263 1886 10309
rect 1858 10235 2846 10263
rect 10210 10235 11198 10263
rect 10210 10189 10238 10235
rect 1474 10161 1694 10189
rect 2914 10161 3134 10189
rect 6754 10161 7358 10189
rect 6754 10115 6782 10161
rect 7330 10152 7358 10161
rect 9826 10161 10238 10189
rect 11170 10189 11198 10235
rect 11170 10161 12062 10189
rect 9826 10152 9854 10161
rect 7330 10124 9854 10152
rect 6562 10087 6782 10115
rect 12034 10115 12062 10161
rect 12034 10087 12254 10115
rect 12706 10087 13118 10115
rect 0 9941 14016 10039
rect 2146 9865 2654 9893
rect 3106 9865 3326 9893
rect 3298 9856 3326 9865
rect 8770 9865 8990 9893
rect 12514 9865 12734 9893
rect 8770 9856 8798 9865
rect 12514 9856 12542 9865
rect 3298 9828 6686 9856
rect 6658 9819 6686 9828
rect 7810 9828 8798 9856
rect 10306 9828 12542 9856
rect 7810 9819 7838 9828
rect 10306 9819 10334 9828
rect 1570 9791 1694 9819
rect 1858 9791 2366 9819
rect 6658 9791 7838 9819
rect 9154 9791 10334 9819
rect 1378 9643 1502 9671
rect 1570 9643 1598 9791
rect 9154 9745 9182 9791
rect 2434 9717 3806 9745
rect 3778 9671 3806 9717
rect 5890 9717 6494 9745
rect 8002 9717 9182 9745
rect 10498 9717 11870 9745
rect 5890 9671 5918 9717
rect 11842 9671 11870 9717
rect 12610 9717 12830 9745
rect 12610 9671 12638 9717
rect 1666 9643 2462 9671
rect 3106 9643 3614 9671
rect 3778 9643 5918 9671
rect 6466 9643 6590 9671
rect 7234 9643 8030 9671
rect 8962 9643 9182 9671
rect 9250 9643 10334 9671
rect 11170 9643 11678 9671
rect 11842 9643 12638 9671
rect 418 9569 1118 9597
rect 418 9449 446 9569
rect 226 9421 446 9449
rect 1090 9449 1118 9569
rect 1474 9523 1502 9643
rect 2434 9597 2462 9643
rect 2265 9569 2352 9597
rect 2434 9569 3038 9597
rect 3490 9523 3518 9597
rect 6658 9569 7166 9597
rect 7257 9569 7344 9597
rect 10114 9569 10238 9597
rect 11458 9569 11582 9597
rect 6658 9560 6686 9569
rect 6082 9532 6686 9560
rect 7618 9532 8222 9560
rect 6082 9523 6110 9532
rect 7618 9523 7646 9532
rect 1474 9495 1982 9523
rect 3394 9495 3518 9523
rect 3778 9495 4478 9523
rect 1954 9486 1982 9495
rect 1954 9458 3230 9486
rect 3202 9449 3230 9458
rect 3778 9449 3806 9495
rect 1090 9421 1310 9449
rect 3202 9421 3806 9449
rect 4450 9449 4478 9495
rect 4834 9495 6110 9523
rect 6946 9495 7646 9523
rect 8194 9523 8222 9532
rect 8194 9495 12734 9523
rect 4834 9449 4862 9495
rect 4450 9421 4862 9449
rect 6178 9421 6782 9449
rect 7714 9421 8126 9449
rect 9346 9421 9566 9449
rect 12825 9421 12912 9449
rect 0 9275 14016 9373
rect 226 9199 446 9227
rect 226 8829 254 9199
rect 418 9079 446 9199
rect 2434 9199 2654 9227
rect 3202 9199 3422 9227
rect 10041 9199 10128 9227
rect 12633 9199 12720 9227
rect 2434 9079 2462 9199
rect 11074 9162 11966 9190
rect 11074 9153 11102 9162
rect 8098 9125 9566 9153
rect 9538 9079 9566 9125
rect 10882 9125 11102 9153
rect 11938 9153 11966 9162
rect 13474 9153 13502 9227
rect 11938 9125 13502 9153
rect 10882 9079 10910 9125
rect 418 9051 2462 9079
rect 2818 9051 2942 9079
rect 6274 9051 6494 9079
rect 9538 9051 10910 9079
rect 11266 9051 11870 9079
rect 2722 8977 2846 9005
rect 2914 8977 2942 9051
rect 11842 9042 11870 9051
rect 12610 9051 13310 9079
rect 13378 9051 13694 9079
rect 13858 9051 13982 9079
rect 12610 9042 12638 9051
rect 11842 9014 12638 9042
rect 3024 8977 3111 9005
rect 3586 8977 3806 9005
rect 3874 8977 4190 9005
rect 6370 8977 7166 9005
rect 7234 8977 7934 9005
rect 8674 8977 9086 9005
rect 11577 8977 11664 9005
rect 12802 8977 12926 9005
rect 2818 8931 2846 8977
rect 12994 8931 13022 9005
rect 2818 8903 3518 8931
rect 3490 8857 3518 8903
rect 4258 8903 6110 8931
rect 8674 8903 9374 8931
rect 11074 8903 11486 8931
rect 4258 8857 4286 8903
rect 3490 8829 4286 8857
rect 11458 8857 11486 8903
rect 12706 8903 13022 8931
rect 12706 8857 12734 8903
rect 11458 8829 12734 8857
rect 13090 8783 13118 9005
rect 6658 8755 7070 8783
rect 7330 8755 7742 8783
rect 8697 8755 8784 8783
rect 12898 8755 13118 8783
rect 13474 8755 13790 8783
rect 0 8609 14016 8707
rect 3010 8533 3902 8561
rect 9922 8533 11102 8561
rect 11458 8533 11774 8561
rect 11746 8524 11774 8533
rect 12802 8533 13022 8561
rect 12802 8524 12830 8533
rect 11746 8496 12830 8524
rect 6082 8459 11582 8487
rect 6082 8413 6110 8459
rect 2050 8385 3518 8413
rect 2050 8339 2078 8385
rect 898 8311 1406 8339
rect 1593 8311 1694 8339
rect 1762 8311 2078 8339
rect 2530 8311 2654 8339
rect 1666 8265 1694 8311
rect 2722 8265 2750 8339
rect 2818 8311 2846 8385
rect 3490 8339 3518 8385
rect 3970 8385 6110 8413
rect 6178 8385 6302 8413
rect 7906 8385 8126 8413
rect 8674 8385 8798 8413
rect 10402 8385 10718 8413
rect 3970 8339 3998 8385
rect 11554 8339 11582 8459
rect 12322 8385 13214 8413
rect 12322 8339 12350 8385
rect 3490 8311 3998 8339
rect 6274 8311 6686 8339
rect 6969 8311 7056 8339
rect 7138 8311 7262 8339
rect 7906 8311 8318 8339
rect 1666 8237 2750 8265
rect 418 8200 1310 8228
rect 418 8191 446 8200
rect 226 8163 446 8191
rect 1282 8191 1310 8200
rect 8674 8191 8702 8339
rect 9346 8191 9374 8339
rect 9442 8311 10238 8339
rect 11074 8311 11486 8339
rect 11554 8311 12350 8339
rect 11458 8265 11486 8311
rect 12418 8265 12446 8339
rect 12514 8311 12638 8339
rect 13186 8311 13214 8385
rect 13282 8265 13310 8339
rect 13378 8311 13502 8339
rect 9922 8237 10142 8265
rect 10617 8237 10704 8265
rect 10809 8237 10896 8265
rect 11458 8237 13310 8265
rect 1282 8163 1502 8191
rect 1954 8163 3326 8191
rect 8674 8163 9086 8191
rect 9346 8163 10814 8191
rect 11650 8163 11870 8191
rect 226 8089 254 8163
rect 1474 8117 1502 8163
rect 11650 8117 11678 8163
rect 322 8089 1406 8117
rect 1474 8089 2462 8117
rect 5913 8089 6000 8117
rect 8194 8089 8414 8117
rect 11170 8089 11678 8117
rect 11746 8089 12062 8117
rect 12144 8089 12231 8117
rect 12322 8089 12734 8117
rect 12898 8089 13598 8117
rect 0 7943 14016 8041
rect 2626 7867 2846 7895
rect 2818 7858 2846 7867
rect 4834 7867 5150 7895
rect 9730 7867 10526 7895
rect 2818 7830 4190 7858
rect 1666 7793 1886 7821
rect 1401 7645 1488 7673
rect 1666 7645 1694 7793
rect 4162 7747 4190 7830
rect 4834 7747 4862 7867
rect 10498 7821 10526 7867
rect 12802 7867 13022 7895
rect 12802 7858 12830 7867
rect 11458 7830 12830 7858
rect 11458 7821 11486 7830
rect 10498 7793 11486 7821
rect 3298 7719 3998 7747
rect 4162 7719 4862 7747
rect 8601 7719 8688 7747
rect 9369 7719 9456 7747
rect 11961 7719 12048 7747
rect 1762 7645 2078 7673
rect 3513 7645 3600 7673
rect 10498 7645 11486 7673
rect 11650 7645 12446 7673
rect 13474 7645 13694 7673
rect 10498 7599 10526 7645
rect 226 7571 1118 7599
rect 8962 7571 10526 7599
rect 11458 7599 11486 7645
rect 11458 7571 13118 7599
rect 13666 7571 13982 7599
rect 226 7451 254 7571
rect 34 7423 254 7451
rect 1090 7451 1118 7571
rect 10594 7497 10814 7525
rect 10786 7488 10814 7497
rect 10786 7460 13406 7488
rect 13378 7451 13406 7460
rect 1090 7423 1310 7451
rect 1954 7423 2558 7451
rect 8578 7423 8798 7451
rect 8866 7423 9566 7451
rect 10617 7423 10704 7451
rect 13378 7423 13598 7451
rect 0 7277 14016 7375
rect 130 7155 158 7229
rect 898 7201 1310 7229
rect 7138 7201 7262 7229
rect 13090 7201 13502 7229
rect 130 7127 350 7155
rect 322 7007 350 7127
rect 2338 7127 4478 7155
rect 7330 7127 10334 7155
rect 2338 7081 2366 7127
rect 7330 7118 7358 7127
rect 6754 7090 7358 7118
rect 1378 7053 2366 7081
rect 5986 7053 6206 7081
rect 1378 7007 1406 7053
rect 6754 7007 6782 7090
rect 9538 7053 9662 7081
rect 322 6979 1406 7007
rect 2530 6979 2654 7007
rect 3010 6979 3518 7007
rect 5122 6979 5630 7007
rect 6178 6979 6782 7007
rect 6873 6979 6960 7007
rect 7042 6979 7454 7007
rect 7714 6979 7838 7007
rect 7906 6979 8414 7007
rect 5122 6933 5150 6979
rect 3874 6905 4190 6933
rect 4930 6905 5150 6933
rect 5602 6933 5630 6979
rect 8482 6933 8510 7007
rect 8592 6979 8679 7007
rect 9154 6979 9662 7007
rect 10329 6979 10416 7007
rect 10512 6979 10599 7007
rect 11362 6979 11678 7007
rect 11746 6979 12158 7007
rect 5602 6905 5822 6933
rect 8482 6905 8894 6933
rect 9250 6905 10238 6933
rect 10210 6896 10238 6905
rect 10690 6905 11294 6933
rect 10690 6896 10718 6905
rect 7234 6868 8318 6896
rect 10210 6868 10718 6896
rect 7234 6859 7262 6868
rect 5602 6831 7262 6859
rect 8290 6859 8318 6868
rect 11266 6859 11294 6905
rect 12226 6905 13406 6933
rect 12226 6859 12254 6905
rect 8290 6831 8990 6859
rect 11266 6831 12254 6859
rect 4546 6794 5246 6822
rect 4546 6785 4574 6794
rect 4354 6757 4574 6785
rect 5218 6785 5246 6794
rect 5218 6757 5438 6785
rect 7330 6757 8222 6785
rect 9922 6757 10142 6785
rect 0 6611 14016 6709
rect 1474 6535 3710 6563
rect 3682 6489 3710 6535
rect 4162 6535 4382 6563
rect 6082 6535 6974 6563
rect 7426 6535 7742 6563
rect 10114 6535 10526 6563
rect 4162 6489 4190 6535
rect 2242 6461 3230 6489
rect 3682 6461 4190 6489
rect 1843 6415 1901 6427
rect 1090 6387 1214 6415
rect 1282 6387 1901 6415
rect 3202 6387 3230 6461
rect 1666 6313 1790 6341
rect 1843 6304 1901 6387
rect 6754 6341 6782 6489
rect 10786 6341 10814 6489
rect 11266 6387 11870 6415
rect 13785 6387 13872 6415
rect 11266 6341 11294 6387
rect 1954 6313 2078 6341
rect 2818 6313 3518 6341
rect 5410 6313 5822 6341
rect 6297 6313 6384 6341
rect 6466 6313 6686 6341
rect 6754 6313 7070 6341
rect 7138 6313 7358 6341
rect 10114 6313 10430 6341
rect 10498 6313 10814 6341
rect 11074 6313 11294 6341
rect 11842 6341 11870 6387
rect 11842 6313 12062 6341
rect 1090 6239 1694 6267
rect 1666 6193 1694 6239
rect 2146 6239 2750 6267
rect 5794 6239 6302 6267
rect 8578 6239 9950 6267
rect 10978 6239 11102 6267
rect 12226 6239 13406 6267
rect 2146 6193 2174 6239
rect 825 6165 912 6193
rect 1666 6165 2174 6193
rect 8578 6119 8606 6239
rect 226 6091 1502 6119
rect 8386 6091 8606 6119
rect 9922 6119 9950 6239
rect 12226 6193 12254 6239
rect 11266 6165 12254 6193
rect 11266 6156 11294 6165
rect 10690 6128 11294 6156
rect 10690 6119 10718 6128
rect 9922 6091 10718 6119
rect 13378 6119 13406 6239
rect 13378 6091 13598 6119
rect 13689 6091 13776 6119
rect 0 5945 14016 6043
rect 1762 5869 2366 5897
rect 6466 5869 6878 5897
rect 7810 5869 9086 5897
rect 12610 5869 12830 5897
rect 13186 5869 13598 5897
rect 9154 5832 10142 5860
rect 2722 5795 5438 5823
rect 5506 5795 7358 5823
rect 8313 5795 8400 5823
rect 5410 5721 5438 5795
rect 6274 5721 6782 5749
rect 7330 5675 7358 5795
rect 9154 5749 9182 5832
rect 10114 5823 10142 5832
rect 12610 5823 12638 5869
rect 10114 5795 12638 5823
rect 7714 5721 8318 5749
rect 8482 5721 9182 5749
rect 3490 5647 3806 5675
rect 4642 5647 5438 5675
rect 6754 5647 7262 5675
rect 7330 5647 7742 5675
rect 9058 5647 9950 5675
rect 11385 5647 11472 5675
rect 11842 5647 12350 5675
rect 1378 5573 3422 5601
rect 3682 5573 4574 5601
rect 6370 5573 6878 5601
rect 7138 5527 7166 5601
rect 4834 5499 6590 5527
rect 6658 5499 7166 5527
rect 7330 5527 7358 5601
rect 7906 5573 8606 5601
rect 7906 5527 7934 5573
rect 7330 5499 7934 5527
rect 8578 5527 8606 5573
rect 9538 5527 9566 5601
rect 10114 5573 11198 5601
rect 8578 5499 9374 5527
rect 9538 5499 9662 5527
rect 6562 5453 6590 5499
rect 9346 5453 9374 5499
rect 10114 5453 10142 5573
rect 11170 5527 11198 5573
rect 12514 5573 13406 5601
rect 12514 5527 12542 5573
rect 11170 5499 12542 5527
rect 5986 5425 6110 5453
rect 6562 5425 8510 5453
rect 9346 5425 10142 5453
rect 13378 5453 13406 5573
rect 13378 5425 13598 5453
rect 0 5279 14016 5377
rect 706 5203 830 5231
rect 1305 5203 1392 5231
rect 9634 5203 9758 5231
rect 7906 5129 8318 5157
rect 8290 5083 8318 5129
rect 8866 5129 9950 5157
rect 8866 5083 8894 5129
rect 3993 5055 4080 5083
rect 8290 5055 8894 5083
rect 10306 5083 10334 5231
rect 10402 5203 10718 5231
rect 12322 5129 12542 5157
rect 12514 5083 12542 5129
rect 10306 5055 10814 5083
rect 12514 5055 12830 5083
rect 12994 5055 13214 5083
rect 825 4981 912 5009
rect 1017 4981 1104 5009
rect 1186 4981 1982 5009
rect 3490 4981 5054 5009
rect 5410 4981 7454 5009
rect 9058 4981 9470 5009
rect 9849 4981 9936 5009
rect 1474 4833 1982 4861
rect 1474 4787 1502 4833
rect 1282 4759 1502 4787
rect 1954 4787 1982 4833
rect 9074 4787 9102 4898
rect 10018 4861 10046 5009
rect 10306 4981 10622 5009
rect 10978 4981 11102 5009
rect 12898 4981 13598 5009
rect 13666 4981 13790 5009
rect 9730 4833 10046 4861
rect 11266 4907 11966 4935
rect 11266 4787 11294 4907
rect 1954 4759 3902 4787
rect 6754 4759 7262 4787
rect 8866 4759 9102 4787
rect 10690 4759 11294 4787
rect 11938 4787 11966 4907
rect 11938 4759 12158 4787
rect 13666 4759 13790 4787
rect 0 4613 14016 4711
rect 825 4537 912 4565
rect 4066 4537 4382 4565
rect 7353 4537 7440 4565
rect 8290 4491 8318 4565
rect 11193 4537 11280 4565
rect 12249 4537 12336 4565
rect 8770 4500 9662 4528
rect 8770 4491 8798 4500
rect 1378 4463 2558 4491
rect 2722 4463 7934 4491
rect 8290 4463 8798 4491
rect 9634 4491 9662 4500
rect 9634 4463 13214 4491
rect 1378 4417 1406 4463
rect 1090 4389 1406 4417
rect 2530 4417 2558 4463
rect 7906 4417 7934 4463
rect 2530 4389 4670 4417
rect 7234 4389 7646 4417
rect 7906 4389 8592 4417
rect 9840 4389 10334 4417
rect 13282 4389 13694 4417
rect 1474 4315 2462 4343
rect 2434 4306 2462 4315
rect 3202 4315 3422 4343
rect 3490 4315 3518 4389
rect 4642 4343 4670 4389
rect 12418 4352 13022 4380
rect 12418 4343 12446 4352
rect 3609 4315 3696 4343
rect 3202 4306 3230 4315
rect 2434 4278 3230 4306
rect 3394 4269 3422 4315
rect 4546 4269 4574 4343
rect 4642 4315 4766 4343
rect 4857 4315 4944 4343
rect 5721 4315 5808 4343
rect 5986 4315 7070 4343
rect 7929 4315 8016 4343
rect 8313 4315 8400 4343
rect 9922 4315 11294 4343
rect 11458 4315 12446 4343
rect 12994 4343 13022 4352
rect 12994 4315 13214 4343
rect 13282 4315 13502 4343
rect 226 4241 926 4269
rect 2169 4241 2256 4269
rect 3394 4241 4574 4269
rect 4738 4269 4766 4315
rect 7522 4276 7646 4304
rect 7522 4269 7550 4276
rect 4738 4241 6686 4269
rect 6777 4241 6864 4269
rect 7426 4241 7550 4269
rect 226 4195 254 4241
rect 34 4167 254 4195
rect 898 4195 926 4241
rect 4546 4195 4574 4241
rect 6658 4195 6686 4241
rect 12514 4195 12542 4269
rect 12706 4241 13118 4269
rect 898 4167 3902 4195
rect 4546 4167 5150 4195
rect 6658 4167 7742 4195
rect 8002 4167 8606 4195
rect 10114 4167 12542 4195
rect 34 4093 62 4167
rect 3874 4121 3902 4167
rect 5122 4158 5150 4167
rect 5122 4130 6494 4158
rect 6466 4121 6494 4130
rect 2914 4093 3230 4121
rect 3298 4093 3806 4121
rect 3874 4093 4958 4121
rect 6466 4093 7454 4121
rect 8002 4093 8030 4167
rect 8578 4093 8606 4167
rect 0 3947 14016 4045
rect 802 3871 1118 3899
rect 1666 3871 2270 3899
rect 5602 3871 5822 3899
rect 6274 3871 6494 3899
rect 9058 3871 9566 3899
rect 9634 3871 10142 3899
rect 10306 3871 10430 3899
rect 9634 3825 9662 3871
rect 10690 3825 10718 3899
rect 10882 3871 11102 3899
rect 12802 3871 13118 3899
rect 13858 3871 13982 3899
rect 7522 3797 8894 3825
rect 9346 3797 9662 3825
rect 10210 3797 10718 3825
rect 12034 3797 12254 3825
rect 7522 3751 7550 3797
rect 1090 3723 1406 3751
rect 2914 3723 3038 3751
rect 3682 3723 7550 3751
rect 8866 3751 8894 3797
rect 12418 3760 13502 3788
rect 12418 3751 12446 3760
rect 8866 3723 12446 3751
rect 13474 3751 13502 3760
rect 13474 3723 13694 3751
rect 13785 3723 13872 3751
rect 1186 3649 1310 3677
rect 1378 3603 1406 3723
rect 1488 3649 1575 3677
rect 2626 3649 3422 3677
rect 7618 3649 7934 3677
rect 8002 3649 8318 3677
rect 8386 3649 9758 3677
rect 8386 3603 8414 3649
rect 1378 3575 1982 3603
rect 7426 3575 8414 3603
rect 8482 3575 9662 3603
rect 8482 3529 8510 3575
rect 9730 3529 9758 3649
rect 9826 3649 9927 3677
rect 10402 3649 10526 3677
rect 9826 3603 9854 3649
rect 10594 3603 10622 3677
rect 9826 3575 10622 3603
rect 10690 3529 10718 3677
rect 11961 3649 12048 3677
rect 12226 3649 12926 3677
rect 12994 3649 13118 3677
rect 13200 3649 13287 3677
rect 12898 3603 12926 3649
rect 12898 3575 13694 3603
rect 4642 3501 6014 3529
rect 7138 3501 8510 3529
rect 9081 3501 9168 3529
rect 9730 3501 10718 3529
rect 10882 3501 12734 3529
rect 4642 3455 4670 3501
rect 4354 3427 4670 3455
rect 5986 3455 6014 3501
rect 10882 3455 10910 3501
rect 5986 3427 6206 3455
rect 6562 3427 10910 3455
rect 12706 3455 12734 3501
rect 12706 3427 13310 3455
rect 0 3281 14016 3379
rect 3682 3205 3902 3233
rect 3874 3159 3902 3205
rect 4354 3205 4574 3233
rect 5698 3205 6014 3233
rect 7042 3205 7262 3233
rect 4354 3159 4382 3205
rect 7234 3196 7262 3205
rect 8002 3205 8222 3233
rect 9154 3205 9374 3233
rect 8002 3196 8030 3205
rect 7234 3168 8030 3196
rect 2914 3131 3518 3159
rect 3874 3131 4382 3159
rect 9346 3159 9374 3205
rect 11650 3205 12062 3233
rect 12418 3205 13022 3233
rect 13113 3205 13200 3233
rect 11650 3196 11678 3205
rect 9922 3168 11678 3196
rect 9922 3159 9950 3168
rect 9346 3131 9950 3159
rect 2914 3085 2942 3131
rect 2242 3057 2942 3085
rect 3490 3085 3518 3131
rect 11842 3094 12542 3122
rect 11842 3085 11870 3094
rect 3490 3057 3710 3085
rect 2242 3011 2270 3057
rect 1474 2983 1886 3011
rect 1968 2983 2055 3011
rect 2169 2983 2270 3011
rect 3010 2983 3518 3011
rect 3682 2937 3710 3057
rect 4642 3057 5630 3085
rect 4642 2937 4670 3057
rect 5602 3011 5630 3057
rect 6082 3057 6686 3085
rect 10690 3057 10910 3085
rect 6082 3011 6110 3057
rect 10882 3011 10910 3057
rect 11650 3057 11870 3085
rect 12514 3085 12542 3094
rect 12514 3057 12734 3085
rect 11650 3011 11678 3057
rect 5602 2983 6110 3011
rect 7234 2983 7934 3011
rect 8002 2983 8414 3011
rect 10114 2983 10334 3011
rect 10882 2983 11678 3011
rect 12130 2983 12638 3011
rect 1666 2909 1886 2937
rect 1858 2900 1886 2909
rect 2338 2909 3422 2937
rect 3682 2909 4670 2937
rect 6658 2909 6878 2937
rect 2338 2900 2366 2909
rect 1858 2872 2366 2900
rect 8002 2863 8030 2983
rect 8578 2909 9086 2937
rect 10498 2909 10622 2937
rect 11842 2909 12062 2937
rect 12153 2909 12240 2937
rect 12322 2909 12542 2937
rect 11842 2863 11870 2909
rect 12322 2863 12350 2909
rect 7042 2835 8510 2863
rect 11842 2835 12350 2863
rect 12610 2863 12638 2983
rect 12706 2937 12734 3057
rect 12898 2983 13310 3011
rect 13378 2983 13886 3011
rect 12706 2909 12830 2937
rect 12898 2863 12926 2983
rect 12610 2835 12926 2863
rect 2242 2761 2462 2789
rect 11074 2761 12830 2789
rect 0 2615 14016 2713
rect 6658 2539 6782 2567
rect 7330 2539 7550 2567
rect 12130 2539 12254 2567
rect 4930 2391 5630 2419
rect 4930 2271 4958 2391
rect 4738 2243 4958 2271
rect 5602 2271 5630 2391
rect 5794 2317 5918 2345
rect 6082 2317 6206 2345
rect 6873 2317 6960 2345
rect 5602 2243 5918 2271
rect 5890 2197 5918 2243
rect 7042 2197 7070 2335
rect 7234 2317 7262 2493
rect 7906 2317 8126 2345
rect 8482 2317 8702 2345
rect 10306 2317 10622 2345
rect 10978 2317 11102 2345
rect 5890 2169 7070 2197
rect 4642 2132 5438 2160
rect 4642 2123 4670 2132
rect 4258 2095 4670 2123
rect 5410 2123 5438 2132
rect 5410 2095 5630 2123
rect 9538 2095 9662 2123
rect 0 1949 14016 2047
rect 2242 1873 2462 1901
rect 2434 1864 2462 1873
rect 3586 1873 3806 1901
rect 4738 1873 4958 1901
rect 3586 1864 3614 1873
rect 2434 1836 3614 1864
rect 4258 1799 4478 1827
rect 2242 1651 3134 1679
rect 4258 1661 4286 1799
rect 4930 1753 4958 1873
rect 8098 1873 8318 1901
rect 9058 1873 9758 1901
rect 8098 1864 8126 1873
rect 5698 1836 8126 1864
rect 5698 1753 5726 1836
rect 8866 1799 9566 1827
rect 4930 1725 5726 1753
rect 9730 1753 9758 1873
rect 13474 1873 13694 1901
rect 11266 1836 12542 1864
rect 11266 1753 11294 1836
rect 12514 1827 12542 1836
rect 13474 1827 13502 1873
rect 12514 1799 13502 1827
rect 9730 1725 11294 1753
rect 4377 1651 4464 1679
rect 5890 1651 8030 1679
rect 11746 1651 12350 1679
rect 1090 1577 2078 1605
rect 2553 1577 2640 1605
rect 3298 1577 3998 1605
rect 1090 1457 1118 1577
rect 2050 1494 2078 1577
rect 3298 1494 3326 1577
rect 2050 1466 3326 1494
rect 898 1429 1118 1457
rect 3970 1457 3998 1577
rect 4564 1457 4592 1633
rect 6201 1577 6288 1605
rect 8290 1577 8414 1605
rect 8578 1577 9566 1605
rect 11458 1577 11966 1605
rect 12898 1577 13310 1605
rect 8578 1494 8606 1577
rect 9538 1531 9566 1577
rect 9538 1503 9950 1531
rect 13570 1503 13790 1531
rect 5890 1466 7262 1494
rect 5890 1457 5918 1466
rect 3970 1429 4190 1457
rect 4354 1429 4592 1457
rect 5122 1429 5918 1457
rect 7234 1457 7262 1466
rect 7618 1466 8606 1494
rect 12322 1466 13022 1494
rect 7618 1457 7646 1466
rect 12322 1457 12350 1466
rect 7234 1429 7646 1457
rect 9657 1429 9744 1457
rect 10594 1429 10718 1457
rect 12130 1429 12350 1457
rect 12994 1457 13022 1466
rect 12994 1429 13214 1457
rect 0 1283 14016 1381
rect 1666 1207 1886 1235
rect 1858 1087 1886 1207
rect 3106 1207 3326 1235
rect 7042 1207 7646 1235
rect 8194 1207 8702 1235
rect 10210 1207 10622 1235
rect 3106 1087 3134 1207
rect 7042 1133 7070 1207
rect 1858 1059 3134 1087
rect 9058 1059 9662 1087
rect 9730 1059 10334 1087
rect 10498 1059 10718 1087
rect 12034 1059 12158 1087
rect 9730 1013 9758 1059
rect 4546 985 5630 1013
rect 5986 985 6110 1013
rect 6658 985 7646 1013
rect 7833 985 7934 1013
rect 8002 985 8990 1013
rect 9250 985 9758 1013
rect 12322 985 12446 1013
rect 7906 939 7934 985
rect 7906 911 9470 939
rect 12706 911 13790 939
rect 7426 800 9566 828
rect 7426 791 7454 800
rect 3874 763 4286 791
rect 7234 763 7454 791
rect 9538 791 9566 800
rect 12706 791 12734 911
rect 9538 763 9758 791
rect 10617 763 10704 791
rect 12514 763 12734 791
rect 13762 791 13790 911
rect 13762 763 13982 791
rect 0 617 14016 715
rect 2626 541 2942 569
rect 4473 541 4560 569
rect 5817 541 5904 569
rect 6274 541 6494 569
rect 6658 541 7358 569
rect 8290 541 8414 569
rect 9058 541 9566 569
rect 10617 541 10704 569
rect 11170 541 11486 569
rect 7330 532 7358 541
rect 7330 504 8030 532
rect 3394 467 4094 495
rect 5506 467 7166 495
rect 3394 421 3422 467
rect 3202 393 3422 421
rect 4066 421 4094 467
rect 8002 421 8030 504
rect 4066 393 6782 421
rect 3106 273 3134 347
rect 3202 319 3230 393
rect 3490 319 3902 347
rect 4066 319 4190 347
rect 4258 319 4286 393
rect 5410 347 5438 393
rect 6754 347 6782 393
rect 4354 273 4382 347
rect 5122 319 5342 347
rect 5410 319 5630 347
rect 5698 319 6686 347
rect 6754 319 6974 347
rect 7042 319 7262 347
rect 5698 273 5726 319
rect 3106 245 5726 273
rect 6946 273 6974 319
rect 7906 273 7934 421
rect 8002 393 9278 421
rect 8578 319 8606 393
rect 8674 273 8702 347
rect 6946 245 8702 273
rect 9250 273 9278 393
rect 9250 245 11006 273
rect 130 171 6878 199
rect 7042 134 8798 162
rect 7042 125 7070 134
rect 3298 97 3518 125
rect 3970 97 4094 125
rect 4930 97 5342 125
rect 6658 97 7070 125
rect 8770 125 8798 134
rect 8770 97 8990 125
rect 0 -49 14016 49
<< metal2 >>
rect 34 7525 62 14652
rect 226 14157 254 14569
rect 226 12973 254 13349
rect 226 11863 254 12251
rect 898 12187 926 12335
rect 802 12159 926 12187
rect 226 11125 254 11743
rect 802 11521 830 12159
rect 1090 11595 1118 14652
rect 1090 11567 1214 11595
rect 802 11493 926 11521
rect 898 11151 926 11493
rect 802 11123 926 11151
rect 226 10027 254 10559
rect 802 10189 830 11123
rect 1186 11077 1214 11567
rect 1090 11049 1214 11077
rect 802 10161 926 10189
rect 898 9819 926 10161
rect 802 9791 926 9819
rect 226 8929 254 9449
rect 802 8857 830 9791
rect 1090 8931 1118 11049
rect 1282 10309 1310 10781
rect 1474 10383 1694 10411
rect 1474 10189 1502 10383
rect 1858 10337 1886 11521
rect 1378 10161 1502 10189
rect 1666 10309 1886 10337
rect 1378 9079 1406 10161
rect 1666 9449 1694 10309
rect 1858 9643 1886 10263
rect 2146 9865 2174 14652
rect 2338 10781 2366 10929
rect 2338 10753 2462 10781
rect 2434 9967 2462 10753
rect 2818 10235 2846 11225
rect 3202 10531 3230 14652
rect 4258 14481 4286 14652
rect 3874 14453 4286 14481
rect 3874 12233 3902 14453
rect 4834 13149 4862 14407
rect 5314 14111 5342 14652
rect 5122 14083 5342 14111
rect 5122 13889 5150 14083
rect 5122 13861 5246 13889
rect 5218 13741 5246 13861
rect 5122 13713 5246 13741
rect 5122 13223 5150 13713
rect 5122 13195 5246 13223
rect 5410 13195 5438 13741
rect 6082 13639 6110 14111
rect 6370 13445 6398 14652
rect 6082 13297 6110 13445
rect 5986 13269 6110 13297
rect 6274 13417 6398 13445
rect 4738 13121 4862 13149
rect 2338 9939 2462 9967
rect 2338 9791 2366 9939
rect 3106 9865 3134 10189
rect 1666 9421 1886 9449
rect 1858 9227 1886 9421
rect 1666 9199 1886 9227
rect 1666 9079 1694 9199
rect 1378 9051 1502 9079
rect 1666 9051 1790 9079
rect 1090 8903 1214 8931
rect 226 8197 254 8857
rect 802 8829 926 8857
rect 898 8191 926 8829
rect 802 8163 926 8191
rect 34 7497 158 7525
rect 34 4781 62 7451
rect 130 7201 158 7497
rect 226 6733 254 8117
rect 322 7155 350 8117
rect 802 7525 830 8163
rect 1186 8117 1214 8903
rect 1090 8089 1214 8117
rect 802 7497 926 7525
rect 898 7201 926 7497
rect 322 7127 542 7155
rect 514 6415 542 7127
rect 226 6387 542 6415
rect 1090 6387 1118 8089
rect 1474 6535 1502 9051
rect 1762 8487 1790 9051
rect 1666 8459 1790 8487
rect 1666 8117 1694 8459
rect 1666 8089 1886 8117
rect 1858 7673 1886 8089
rect 1762 7645 1886 7673
rect 1762 6859 1790 7645
rect 1762 6831 1886 6859
rect 226 6245 254 6387
rect 226 5823 254 6119
rect 226 5795 350 5823
rect 322 4861 350 5795
rect 226 4833 350 4861
rect 226 4195 254 4833
rect 226 4167 350 4195
rect 34 389 62 4121
rect 322 3677 350 4167
rect 226 3649 350 3677
rect 226 3439 254 3649
rect 706 3233 734 5231
rect 898 4537 926 6193
rect 1282 5601 1310 6415
rect 1858 6387 1886 6831
rect 1762 5869 1790 6341
rect 2050 6193 2078 8339
rect 1954 6165 2078 6193
rect 1090 5573 1310 5601
rect 322 3205 734 3233
rect 322 2567 350 3205
rect 226 2539 350 2567
rect 226 2341 254 2539
rect 802 1383 830 3899
rect 1090 3723 1118 5573
rect 1378 5203 1406 5601
rect 1282 3649 1310 4787
rect 1474 2983 1502 5009
rect 1954 4981 1982 6165
rect 2338 5869 2366 9597
rect 2818 8783 2846 9079
rect 2722 8755 2846 8783
rect 3010 8783 3038 9597
rect 3394 9199 3422 9523
rect 3010 8755 3134 8783
rect 2626 7867 2654 8339
rect 2722 8311 2750 8755
rect 3106 8385 3134 8755
rect 3298 7719 3326 8191
rect 3586 7451 3614 11003
rect 4738 10929 4766 13121
rect 4738 10901 4862 10929
rect 4834 10753 4862 10901
rect 3874 8533 3902 9005
rect 5026 7867 5054 13075
rect 5218 13047 5246 13195
rect 5986 12483 6014 13269
rect 5986 12455 6110 12483
rect 6082 12307 6110 12455
rect 5218 11447 5246 11669
rect 5122 11419 5246 11447
rect 5410 11447 5438 12261
rect 5410 11419 5534 11447
rect 5122 11197 5150 11419
rect 5506 10531 5534 11419
rect 5794 10901 5822 11447
rect 6178 8385 6206 9449
rect 6274 9051 6302 13417
rect 6850 11863 6878 13001
rect 7522 12853 7550 14652
rect 8578 14379 8606 14652
rect 8386 13075 8414 14185
rect 7234 12825 7550 12853
rect 8290 13047 8414 13075
rect 7234 12261 7262 12825
rect 7522 12307 7550 12779
rect 7234 12233 7358 12261
rect 6562 11197 6590 11669
rect 6562 9643 6590 10115
rect 6850 9495 6974 9523
rect 2530 6979 2558 7451
rect 3490 7423 3614 7451
rect 2722 5795 2750 6267
rect 2242 3871 2270 4269
rect 2914 3723 2942 4121
rect 1954 2983 1982 3603
rect 2242 2863 2270 3011
rect 2146 2835 2270 2863
rect 2146 2049 2174 2835
rect 2146 2021 2270 2049
rect 2242 1873 2270 2021
rect 2434 1679 2462 2789
rect 2338 1651 2462 1679
rect 3106 1651 3134 3011
rect 3298 2863 3326 4121
rect 3490 3677 3518 7423
rect 5986 7053 6014 8117
rect 6658 7821 6686 8783
rect 6562 7793 6686 7821
rect 3682 4713 3710 5601
rect 3874 4759 3902 6933
rect 3682 4685 3902 4713
rect 3394 3649 3518 3677
rect 3490 2983 3518 3649
rect 3682 3205 3710 4343
rect 3874 3825 3902 4685
rect 4066 4537 4094 5083
rect 3874 3797 3998 3825
rect 3970 3159 3998 3797
rect 4642 3751 4670 4343
rect 4930 4315 4958 6933
rect 6562 6859 6590 7793
rect 6850 7081 6878 9495
rect 7042 8311 7070 12113
rect 7330 9569 7358 12233
rect 7714 11641 7742 12113
rect 8290 12039 8318 13047
rect 8290 12011 8414 12039
rect 8386 11863 8414 12011
rect 8578 11743 8606 13001
rect 9058 11891 9086 13075
rect 9634 12557 9662 14652
rect 10690 12631 10718 14652
rect 11746 13149 11774 14652
rect 11650 13121 11774 13149
rect 12802 13001 12830 14652
rect 13954 14333 13982 14652
rect 13474 14305 13982 14333
rect 12706 12973 12830 13001
rect 9538 12529 9662 12557
rect 10594 12603 10718 12631
rect 10594 12039 10622 12603
rect 10594 12011 10718 12039
rect 8482 11715 8606 11743
rect 8770 11863 9086 11891
rect 10690 11863 10718 12011
rect 7618 10309 7646 11003
rect 8002 10383 8030 11447
rect 8194 10975 8222 11447
rect 8482 11151 8510 11715
rect 8770 11197 8798 11863
rect 8482 11123 8606 11151
rect 9250 11123 9278 11743
rect 10882 11669 10910 12557
rect 12706 12529 12734 12739
rect 12994 12409 13022 13349
rect 12898 12381 13022 12409
rect 12898 11669 12926 12381
rect 10786 11641 10910 11669
rect 12802 11641 12926 11669
rect 8578 10531 8606 11123
rect 9442 10383 9470 11447
rect 9634 11299 9662 11447
rect 9634 11271 9758 11299
rect 9730 10337 9758 11271
rect 10786 11003 10814 11641
rect 10786 10975 10910 11003
rect 10690 10707 10718 10855
rect 9634 10309 9758 10337
rect 10594 10679 10718 10707
rect 8962 9643 8990 9893
rect 7330 8413 7358 8783
rect 7330 8385 7454 8413
rect 8098 8385 8126 9449
rect 8770 8385 8798 8783
rect 7234 8191 7262 8339
rect 7138 8163 7262 8191
rect 7138 7377 7166 8163
rect 7426 7525 7454 8385
rect 7330 7497 7454 7525
rect 7138 7349 7262 7377
rect 7234 7201 7262 7349
rect 7330 7155 7358 7497
rect 6802 7053 6878 7081
rect 7138 7127 7358 7155
rect 5410 6313 5438 6785
rect 5602 4417 5630 6859
rect 6562 6831 6686 6859
rect 6370 6313 6494 6341
rect 6658 6313 6686 6831
rect 6802 6489 6830 7053
rect 6946 6535 6974 7007
rect 6802 6461 6878 6489
rect 5506 4389 5630 4417
rect 5506 3825 5534 4389
rect 5794 3871 5822 4343
rect 5506 3797 5630 3825
rect 4642 3723 4766 3751
rect 3874 3131 3998 3159
rect 3298 2835 3422 2863
rect 226 1355 830 1383
rect 226 1243 254 1355
rect 130 0 158 199
rect 898 0 926 1457
rect 1666 0 1694 1235
rect 2338 495 2366 1651
rect 3394 1605 3422 2835
rect 2626 541 2654 1605
rect 3298 1577 3422 1605
rect 3298 1207 3326 1577
rect 2338 467 2462 495
rect 2434 0 2462 467
rect 3874 319 3902 3131
rect 4258 1235 4286 2123
rect 4450 1799 4478 3455
rect 4738 1679 4766 3723
rect 5602 2095 5630 3797
rect 5986 2419 6014 5453
rect 6274 3871 6302 6267
rect 6466 5869 6494 6313
rect 6850 5573 6878 6461
rect 7138 6267 7166 7127
rect 7330 6313 7358 6785
rect 7714 6535 7742 7007
rect 8386 6979 8414 8117
rect 8674 7599 8702 7747
rect 8674 7571 8750 7599
rect 8578 6979 8606 7451
rect 8722 6933 8750 7571
rect 9058 7525 9086 9005
rect 9346 8903 9374 9449
rect 9442 7599 9470 7747
rect 9634 7673 9662 10309
rect 10114 8783 10142 9597
rect 9922 8755 10142 8783
rect 9922 8533 9950 8755
rect 10594 8561 10622 10679
rect 10594 8533 10718 8561
rect 10690 8385 10718 8533
rect 9346 7571 9470 7599
rect 9538 7645 9662 7673
rect 9058 7497 9182 7525
rect 8674 6905 8750 6933
rect 8866 6905 8894 7451
rect 7138 6239 7262 6267
rect 6658 3825 6686 5527
rect 6562 3797 6686 3825
rect 6562 3233 6590 3797
rect 6562 3205 6686 3233
rect 6658 3057 6686 3205
rect 6658 2539 6686 2937
rect 5986 2391 6590 2419
rect 5890 1975 5918 2345
rect 4450 1651 4766 1679
rect 4162 1207 4286 1235
rect 4162 319 4190 1207
rect 4354 319 4382 1457
rect 4738 1087 4766 1651
rect 5794 1947 5918 1975
rect 4738 1059 4862 1087
rect 4546 541 4574 1013
rect 4834 569 4862 1059
rect 4738 541 4862 569
rect 4738 393 4766 541
rect 5122 319 5150 1457
rect 5794 939 5822 1947
rect 6082 985 6110 2345
rect 5794 911 5918 939
rect 5890 541 5918 911
rect 6274 541 6302 1605
rect 6562 1531 6590 2391
rect 6562 1503 6686 1531
rect 6658 985 6686 1503
rect 3202 97 3326 125
rect 3970 97 4094 125
rect 4738 97 4958 125
rect 3202 0 3230 97
rect 3970 0 3998 97
rect 4738 0 4766 97
rect 5506 0 5534 495
rect 6658 319 6686 569
rect 6850 171 6878 4269
rect 7042 3205 7070 4343
rect 7234 4269 7262 6239
rect 8386 5795 8414 6119
rect 7426 4537 7454 5009
rect 7618 4537 8030 4565
rect 7618 4389 7646 4537
rect 7234 4241 7310 4269
rect 7138 3501 7166 4195
rect 7282 3455 7310 4241
rect 7234 3427 7310 3455
rect 7042 2345 7070 2863
rect 7234 2465 7262 3427
rect 7426 2835 7454 4269
rect 7714 4167 7742 4343
rect 6946 2317 7070 2345
rect 6274 97 6686 125
rect 6274 0 6302 97
rect 7042 0 7070 1161
rect 7234 319 7262 791
rect 7522 569 7550 2567
rect 7906 1651 7934 4417
rect 8098 4343 8126 5157
rect 8290 4537 8318 5749
rect 8482 5425 8510 5749
rect 8002 4315 8126 4343
rect 8386 4315 8414 4565
rect 8290 2789 8318 3677
rect 8194 2761 8318 2789
rect 8194 2049 8222 2761
rect 8482 2715 8510 2863
rect 8434 2687 8510 2715
rect 8194 2021 8318 2049
rect 8290 1873 8318 2021
rect 8290 1457 8318 1605
rect 8194 1429 8318 1457
rect 7522 541 7838 569
rect 7810 0 7838 541
rect 7906 393 7934 1013
rect 8194 717 8222 1429
rect 8434 1161 8462 2687
rect 8434 1133 8510 1161
rect 8194 689 8318 717
rect 8290 541 8318 689
rect 8482 393 8510 1133
rect 8578 1087 8606 4121
rect 8674 3825 8702 6905
rect 9154 6859 9182 7497
rect 9346 7007 9374 7571
rect 9538 7053 9566 7645
rect 9346 6979 9470 7007
rect 9058 6831 9182 6859
rect 9058 5869 9086 6831
rect 8866 4343 8894 4787
rect 9058 4389 9086 5675
rect 8866 4315 9086 4343
rect 9058 3871 9086 4315
rect 9442 3973 9470 6979
rect 9922 6859 9950 8265
rect 10402 7497 10622 7525
rect 10402 6979 10430 7497
rect 10690 7081 10718 8265
rect 10882 8237 10910 10975
rect 11074 10485 11102 11595
rect 12706 10827 12734 10909
rect 11074 10457 11198 10485
rect 11170 9523 11198 10457
rect 11074 9495 11198 9523
rect 11074 8311 11102 9495
rect 11458 8533 11486 9597
rect 10690 7053 10814 7081
rect 9826 6831 9950 6859
rect 9826 6267 9854 6831
rect 10114 6313 10142 6785
rect 10498 6535 10526 7007
rect 10786 6415 10814 7053
rect 10690 6387 10814 6415
rect 9826 6239 9950 6267
rect 9634 5203 9662 5527
rect 9922 5129 9950 6239
rect 9442 3945 9566 3973
rect 8674 3797 8798 3825
rect 8770 3677 8798 3797
rect 8770 3649 8894 3677
rect 8866 3085 8894 3649
rect 9154 3205 9182 3529
rect 8770 3057 8894 3085
rect 8770 2863 8798 3057
rect 8674 2835 8798 2863
rect 8674 2567 8702 2835
rect 8674 2539 8894 2567
rect 8674 2197 8702 2345
rect 8674 2169 8750 2197
rect 8722 1531 8750 2169
rect 8866 1799 8894 2539
rect 8674 1503 8750 1531
rect 8674 1207 8702 1503
rect 8578 1059 8798 1087
rect 9058 1059 9086 2937
rect 8770 347 8798 1059
rect 8578 319 8798 347
rect 8578 0 8606 319
rect 9346 0 9374 3825
rect 9538 3455 9566 3945
rect 9730 3677 9758 4861
rect 9922 4565 9950 5009
rect 9922 4537 10142 4565
rect 9634 3649 9854 3677
rect 9634 3575 9662 3649
rect 9538 3427 9662 3455
rect 9634 2271 9662 3427
rect 9538 2243 9662 2271
rect 9538 541 9566 2243
rect 9922 1503 9950 4343
rect 10114 3501 10142 4537
rect 10306 2317 10334 5297
rect 10402 1827 10430 3899
rect 10498 3649 10526 6119
rect 10690 5203 10718 6387
rect 10978 5157 11006 6267
rect 11458 5453 11486 5675
rect 11650 5453 11678 9671
rect 12322 8561 12350 10411
rect 12706 9865 12734 10115
rect 12802 9717 12830 11641
rect 12994 10485 13022 11519
rect 13186 10633 13214 13959
rect 13186 10605 13310 10633
rect 12994 10457 13214 10485
rect 12898 10263 12926 10411
rect 12898 10235 13022 10263
rect 12994 9671 13022 10235
rect 12898 9643 13022 9671
rect 12706 9495 12734 9567
rect 12322 8533 12542 8561
rect 12514 8311 12542 8533
rect 12706 8191 12734 9227
rect 12898 8977 12926 9643
rect 12898 8385 12926 8783
rect 11074 5425 11678 5453
rect 11074 5269 11102 5425
rect 10978 5129 11294 5157
rect 10786 5055 10910 5083
rect 10690 3871 10718 4787
rect 10882 3751 10910 5055
rect 11074 3871 11102 5009
rect 11266 4537 11294 5129
rect 10882 3723 11006 3751
rect 10690 3057 10718 3529
rect 10978 3011 11006 3723
rect 10882 2983 11006 3011
rect 10306 1799 10430 1827
rect 9730 763 9758 1457
rect 10306 1161 10334 1799
rect 10594 1207 10622 2937
rect 10306 1133 10430 1161
rect 10402 569 10430 1133
rect 10690 1059 10718 1457
rect 10882 1161 10910 2983
rect 11074 2317 11102 2789
rect 11650 2567 11678 5425
rect 11842 3011 11870 8191
rect 12610 8163 12734 8191
rect 12034 7719 12062 8117
rect 12130 6979 12158 8117
rect 12034 3797 12062 6341
rect 12322 5749 12350 8117
rect 12610 7525 12638 8163
rect 12898 7525 12926 8117
rect 12994 7867 13022 8957
rect 13186 8487 13214 10457
rect 13282 10383 13310 10605
rect 13474 10531 13502 14305
rect 13762 12101 13886 12129
rect 13858 11891 13886 12101
rect 13762 11863 13886 11891
rect 13762 10781 13790 11863
rect 13762 10753 13886 10781
rect 13858 10559 13886 10753
rect 13762 10531 13886 10559
rect 13570 10115 13598 10299
rect 13474 10087 13598 10115
rect 13474 9199 13502 10087
rect 13762 9523 13790 10531
rect 13762 9495 13886 9523
rect 13186 8459 13262 8487
rect 13090 7571 13118 8347
rect 13234 7525 13262 8459
rect 13378 7599 13406 9079
rect 13474 7645 13502 8783
rect 13378 7571 13502 7599
rect 12610 7497 12734 7525
rect 12898 7497 13022 7525
rect 12226 5721 12350 5749
rect 12226 4491 12254 5721
rect 12322 5527 12350 5675
rect 12322 5499 12446 5527
rect 12418 4861 12446 5499
rect 12322 4833 12446 4861
rect 12322 4537 12350 4833
rect 12226 4463 12350 4491
rect 12034 3011 12062 3677
rect 12322 3085 12350 4463
rect 12706 4417 12734 7497
rect 12802 5833 12830 5907
rect 12610 4389 12734 4417
rect 12610 3677 12638 4389
rect 12994 4343 13022 7497
rect 13186 7497 13262 7525
rect 13186 5055 13214 7497
rect 13474 7201 13502 7571
rect 13378 6905 13406 7127
rect 13666 6785 13694 7737
rect 13858 7673 13886 9495
rect 13954 9051 13982 14203
rect 13810 7645 13886 7673
rect 13810 6859 13838 7645
rect 13810 6831 13886 6859
rect 13378 6757 13694 6785
rect 13378 5009 13406 6757
rect 13570 5869 13598 6517
rect 13858 6387 13886 6831
rect 13570 5269 13598 5453
rect 12898 4315 13022 4343
rect 13186 4981 13406 5009
rect 13762 4981 13790 6119
rect 13186 4315 13214 4981
rect 13666 4389 13694 4787
rect 12898 3751 12926 4315
rect 13090 3871 13118 4269
rect 12898 3723 13118 3751
rect 12610 3649 12734 3677
rect 12322 3057 12446 3085
rect 11842 2983 11966 3011
rect 12034 2983 12158 3011
rect 11650 2539 11774 2567
rect 11746 1651 11774 2539
rect 11938 1605 11966 2983
rect 12226 2539 12254 2937
rect 12418 2493 12446 3057
rect 12322 2465 12446 2493
rect 12322 1901 12350 2465
rect 12322 1873 12542 1901
rect 10882 1133 11006 1161
rect 10114 541 10430 569
rect 10690 541 10718 791
rect 10114 0 10142 541
rect 10978 495 11006 1133
rect 11458 541 11486 1605
rect 11746 1577 11966 1605
rect 11746 495 11774 1577
rect 12130 1059 12158 1457
rect 12322 985 12350 1679
rect 12514 763 12542 1873
rect 12706 1457 12734 3649
rect 12994 3205 13022 3677
rect 13090 3159 13118 3723
rect 13186 3205 13214 3677
rect 13282 3427 13310 3955
rect 13090 3131 13214 3159
rect 12802 2909 12926 2937
rect 12898 1577 12926 2909
rect 12706 1429 12830 1457
rect 12802 569 12830 1429
rect 10882 467 11006 495
rect 11650 467 11774 495
rect 12418 541 12830 569
rect 10882 0 10910 467
rect 11650 0 11678 467
rect 12418 0 12446 541
rect 13186 0 13214 3131
rect 13474 877 13502 4343
rect 13762 3751 13790 4565
rect 13954 3871 13982 7599
rect 13762 3723 13886 3751
rect 13666 3317 13694 3603
rect 13858 2271 13886 3011
rect 13858 2243 13982 2271
rect 13666 1873 13694 2125
rect 13762 1452 13790 1531
rect 13954 1383 13982 2243
rect 13858 1355 13982 1383
rect 13858 717 13886 1355
rect 13762 689 13886 717
rect 13762 267 13790 689
rect 13954 0 13982 791
<< metal3 >>
rect 0 14525 270 14585
rect 0 13305 270 13365
rect 0 12207 270 12267
rect 0 11109 270 11169
rect 0 10011 270 10071
rect 0 8913 270 8973
rect 210 7875 270 8241
rect 0 7815 270 7875
rect 0 6717 270 6777
rect 210 5679 270 6289
rect 0 5619 270 5679
rect 18 4581 78 4825
rect 0 4521 160 4581
rect 0 3423 270 3483
rect 0 2325 270 2385
rect 0 1227 270 1287
rect 18 189 78 433
rect 0 129 160 189
rect 400 0 600 14652
rect 1600 0 1800 14652
rect 2800 0 3000 14652
rect 4000 0 4200 14652
rect 5200 0 5400 14652
rect 6400 0 6600 14652
rect 7600 0 7800 14652
rect 7986 4521 8430 4581
rect 8800 0 9000 14652
rect 10000 0 10200 14652
rect 10290 5253 11118 5313
rect 11200 0 11400 14652
rect 12400 0 12600 14652
rect 13856 14525 14016 14585
rect 13600 14095 13800 14405
rect 13938 14159 13998 14525
rect 13170 13915 14016 13975
rect 13600 13485 13800 13795
rect 12978 13305 14016 13365
rect 13600 12875 13800 13185
rect 12690 12695 14016 12755
rect 13600 12265 13800 12575
rect 13746 12085 14016 12145
rect 13600 11655 13800 11965
rect 12978 11475 14016 11535
rect 13600 11045 13800 11355
rect 12690 10865 14016 10925
rect 13600 10435 13800 10745
rect 13554 10255 14016 10315
rect 13600 9703 13800 10135
rect 12690 9523 14016 9583
rect 13600 9093 13800 9403
rect 12978 8913 14016 8973
rect 13600 8483 13800 8793
rect 13074 8303 14016 8363
rect 13600 7873 13800 8183
rect 13650 7693 14016 7753
rect 13600 7263 13800 7573
rect 13362 7083 14016 7143
rect 13600 6653 13800 6963
rect 13554 6473 14016 6533
rect 13600 6043 13800 6353
rect 12786 5863 14016 5923
rect 13600 5433 13800 5743
rect 13554 5253 14016 5313
rect 13600 4701 13800 5133
rect 13746 4521 14016 4581
rect 13600 4091 13800 4401
rect 13266 3911 14016 3971
rect 13600 3481 13800 3791
rect 13650 3301 14016 3361
rect 13600 2871 13800 3181
rect 12882 2691 14016 2751
rect 13600 2261 13800 2571
rect 13650 2081 14016 2141
rect 13600 1651 13800 1961
rect 13746 1471 14016 1531
rect 13600 1041 13800 1351
rect 13458 861 14016 921
rect 13600 431 13800 741
rect 13746 251 14016 311
use M2M3_PR  M2M3_PR_68
timestamp 1626908933
transform 1 0 48 0 1 403
box -33 -37 33 37
use M2M3_PR  M2M3_PR_26
timestamp 1626908933
transform 1 0 48 0 1 403
box -33 -37 33 37
use M1M2_PR  M1M2_PR_929
timestamp 1626908933
transform 1 0 144 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_464
timestamp 1626908933
transform 1 0 144 0 1 185
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_254
timestamp 1626908933
transform 1 0 192 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_251
timestamp 1626908933
transform 1 0 0 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_84
timestamp 1626908933
transform 1 0 192 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_81
timestamp 1626908933
transform 1 0 0 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_163
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_81
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_149
timestamp 1626908933
transform 1 0 0 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_36
timestamp 1626908933
transform 1 0 0 0 1 0
box -38 -49 230 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_65
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_184
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_65
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_184
timestamp 1626908933
transform 1 0 500 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_92
timestamp 1626908933
transform 1 0 768 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_102
timestamp 1626908933
transform 1 0 96 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_195
timestamp 1626908933
transform 1 0 768 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_205
timestamp 1626908933
transform 1 0 96 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_119
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_239
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_250
timestamp 1626908933
transform 1 0 1248 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_80
timestamp 1626908933
transform 1 0 1248 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_148
timestamp 1626908933
transform 1 0 1536 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_35
timestamp 1626908933
transform 1 0 1536 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_230
timestamp 1626908933
transform 1 0 864 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_110
timestamp 1626908933
transform 1 0 864 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_185
timestamp 1626908933
transform 1 0 1344 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_82
timestamp 1626908933
transform 1 0 1344 0 -1 1332
box -38 -49 806 715
use prbs_generator_syn_VIA3  prbs_generator_syn_VIA3_1
timestamp 1626908933
transform 1 0 1761 0 1 23
box -39 -26 39 26
use prbs_generator_syn_VIA3  prbs_generator_syn_VIA3_0
timestamp 1626908933
transform 1 0 1761 0 1 23
box -39 -26 39 26
use prbs_generator_syn_VIA2  prbs_generator_syn_VIA2_1
timestamp 1626908933
transform 1 0 1761 0 1 16
box -39 -33 39 33
use prbs_generator_syn_VIA2  prbs_generator_syn_VIA2_0
timestamp 1626908933
transform 1 0 1761 0 1 16
box -39 -33 39 33
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_180
timestamp 1626908933
transform 1 0 1728 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_77
timestamp 1626908933
transform 1 0 1728 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_162
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_157
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_80
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_75
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_173
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_54
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_173
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_54
timestamp 1626908933
transform 1 0 2900 0 1 666
box -100 -49 100 49
use M1M2_PR  M1M2_PR_708
timestamp 1626908933
transform 1 0 2640 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_243
timestamp 1626908933
transform 1 0 2640 0 1 555
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_255
timestamp 1626908933
transform 1 0 2784 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_85
timestamp 1626908933
transform 1 0 2784 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_150
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_37
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_71
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_174
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_95
timestamp 1626908933
transform 1 0 2112 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_215
timestamp 1626908933
transform 1 0 2112 0 -1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_878
timestamp 1626908933
transform 1 0 3312 0 1 111
box -32 -32 32 32
use M1M2_PR  M1M2_PR_413
timestamp 1626908933
transform 1 0 3312 0 1 111
box -32 -32 32 32
use L1M1_PR  L1M1_PR_957
timestamp 1626908933
transform 1 0 3504 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_455
timestamp 1626908933
transform 1 0 3504 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_992
timestamp 1626908933
transform 1 0 3120 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_490
timestamp 1626908933
transform 1 0 3120 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_761
timestamp 1626908933
transform 1 0 3216 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_259
timestamp 1626908933
transform 1 0 3216 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_589
timestamp 1626908933
transform 1 0 3504 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_87
timestamp 1626908933
transform 1 0 3504 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_294
timestamp 1626908933
transform 1 0 2928 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_796
timestamp 1626908933
transform 1 0 2928 0 1 555
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_62
timestamp 1626908933
transform 1 0 3360 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_165
timestamp 1626908933
transform 1 0 3360 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_78
timestamp 1626908933
transform 1 0 3552 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_198
timestamp 1626908933
transform 1 0 3552 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_3
timestamp 1626908933
transform -1 0 3552 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_35
timestamp 1626908933
transform -1 0 3552 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_36
timestamp 1626908933
transform 1 0 3936 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_4
timestamp 1626908933
transform 1 0 3936 0 1 0
box -38 -49 710 715
use L1M1_PR  L1M1_PR_956
timestamp 1626908933
transform 1 0 3984 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_454
timestamp 1626908933
transform 1 0 3984 0 1 111
box -29 -23 29 23
use M1M2_PR  M1M2_PR_555
timestamp 1626908933
transform 1 0 3888 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_90
timestamp 1626908933
transform 1 0 3888 0 1 333
box -32 -32 32 32
use prbs_generator_syn_VIA7  prbs_generator_syn_VIA7_3
timestamp 1626908933
transform 1 0 4113 0 1 23
box -87 -26 87 26
use prbs_generator_syn_VIA7  prbs_generator_syn_VIA7_1
timestamp 1626908933
transform 1 0 4113 0 1 23
box -87 -26 87 26
use prbs_generator_syn_VIA6  prbs_generator_syn_VIA6_3
timestamp 1626908933
transform 1 0 4113 0 1 16
box -87 -33 87 33
use prbs_generator_syn_VIA6  prbs_generator_syn_VIA6_1
timestamp 1626908933
transform 1 0 4113 0 1 16
box -87 -33 87 33
use M1M2_PR  M1M2_PR_877
timestamp 1626908933
transform 1 0 4080 0 1 111
box -32 -32 32 32
use M1M2_PR  M1M2_PR_412
timestamp 1626908933
transform 1 0 4080 0 1 111
box -32 -32 32 32
use L1M1_PR  L1M1_PR_586
timestamp 1626908933
transform 1 0 4080 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_84
timestamp 1626908933
transform 1 0 4080 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_759
timestamp 1626908933
transform 1 0 4272 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_257
timestamp 1626908933
transform 1 0 4272 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_553
timestamp 1626908933
transform 1 0 4176 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_88
timestamp 1626908933
transform 1 0 4176 0 1 333
box -32 -32 32 32
use L1M1_PR  L1M1_PR_990
timestamp 1626908933
transform 1 0 4368 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_488
timestamp 1626908933
transform 1 0 4368 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_911
timestamp 1626908933
transform 1 0 4368 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_446
timestamp 1626908933
transform 1 0 4368 0 1 333
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_70
timestamp 1626908933
transform 1 0 4608 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_190
timestamp 1626908933
transform 1 0 4608 0 1 0
box -38 -49 422 715
use M1M2_PR  M1M2_PR_203
timestamp 1626908933
transform 1 0 4752 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_245
timestamp 1626908933
transform 1 0 4560 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_668
timestamp 1626908933
transform 1 0 4752 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_710
timestamp 1626908933
transform 1 0 4560 0 1 555
box -32 -32 32 32
use L1M1_PR  L1M1_PR_297
timestamp 1626908933
transform 1 0 4560 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_799
timestamp 1626908933
transform 1 0 4560 0 1 555
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_79
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_161
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use M1M2_PR  M1M2_PR_411
timestamp 1626908933
transform 1 0 4944 0 1 111
box -32 -32 32 32
use M1M2_PR  M1M2_PR_876
timestamp 1626908933
transform 1 0 4944 0 1 111
box -32 -32 32 32
use L1M1_PR  L1M1_PR_955
timestamp 1626908933
transform 1 0 5328 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_583
timestamp 1626908933
transform 1 0 5328 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_453
timestamp 1626908933
transform 1 0 5328 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_81
timestamp 1626908933
transform 1 0 5328 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_549
timestamp 1626908933
transform 1 0 5136 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_84
timestamp 1626908933
transform 1 0 5136 0 1 333
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_162
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_43
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_162
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_43
timestamp 1626908933
transform 1 0 5300 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_151
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_38
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 230 715
use L1M1_PR  L1M1_PR_755
timestamp 1626908933
transform 1 0 5616 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_253
timestamp 1626908933
transform 1 0 5616 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_875
timestamp 1626908933
transform 1 0 5520 0 1 481
box -32 -32 32 32
use M1M2_PR  M1M2_PR_410
timestamp 1626908933
transform 1 0 5520 0 1 481
box -32 -32 32 32
use L1M1_PR  L1M1_PR_986
timestamp 1626908933
transform 1 0 5712 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_484
timestamp 1626908933
transform 1 0 5712 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_800
timestamp 1626908933
transform 1 0 5904 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_298
timestamp 1626908933
transform 1 0 5904 0 1 555
box -29 -23 29 23
use M1M2_PR  M1M2_PR_712
timestamp 1626908933
transform 1 0 5904 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_247
timestamp 1626908933
transform 1 0 5904 0 1 555
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_253
timestamp 1626908933
transform 1 0 5952 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_83
timestamp 1626908933
transform 1 0 5952 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_5
timestamp 1626908933
transform 1 0 5280 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_37
timestamp 1626908933
transform 1 0 5280 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_37
timestamp 1626908933
transform -1 0 6048 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_0
timestamp 1626908933
transform -1 0 6048 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_33
timestamp 1626908933
transform 1 0 6048 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_146
timestamp 1626908933
transform 1 0 6048 0 -1 1332
box -38 -49 230 715
use M1M2_PR  M1M2_PR_249
timestamp 1626908933
transform 1 0 6288 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_714
timestamp 1626908933
transform 1 0 6288 0 1 555
box -32 -32 32 32
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_15
timestamp 1626908933
transform 1 0 6500 0 1 23
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_7
timestamp 1626908933
transform 1 0 6500 0 1 23
box -100 -26 100 26
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_15
timestamp 1626908933
transform 1 0 6500 0 1 16
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_7
timestamp 1626908933
transform 1 0 6500 0 1 16
box -100 -33 100 33
use M1M2_PR  M1M2_PR_874
timestamp 1626908933
transform 1 0 6672 0 1 111
box -32 -32 32 32
use M1M2_PR  M1M2_PR_409
timestamp 1626908933
transform 1 0 6672 0 1 111
box -32 -32 32 32
use L1M1_PR  L1M1_PR_985
timestamp 1626908933
transform 1 0 6672 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_753
timestamp 1626908933
transform 1 0 6768 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_483
timestamp 1626908933
transform 1 0 6672 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_251
timestamp 1626908933
transform 1 0 6768 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_907
timestamp 1626908933
transform 1 0 6672 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_442
timestamp 1626908933
transform 1 0 6672 0 1 333
box -32 -32 32 32
use L1M1_PR  L1M1_PR_802
timestamp 1626908933
transform 1 0 6480 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_300
timestamp 1626908933
transform 1 0 6480 0 1 555
box -29 -23 29 23
use M1M2_PR  M1M2_PR_906
timestamp 1626908933
transform 1 0 6672 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_441
timestamp 1626908933
transform 1 0 6672 0 1 555
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_44
timestamp 1626908933
transform 1 0 6240 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_147
timestamp 1626908933
transform 1 0 6240 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_64
timestamp 1626908933
transform 1 0 6048 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_184
timestamp 1626908933
transform 1 0 6048 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_6
timestamp 1626908933
transform -1 0 7104 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_38
timestamp 1626908933
transform -1 0 7104 0 1 0
box -38 -49 710 715
use M1M2_PR  M1M2_PR_928
timestamp 1626908933
transform 1 0 6864 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_463
timestamp 1626908933
transform 1 0 6864 0 1 185
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_249
timestamp 1626908933
transform 1 0 7008 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_79
timestamp 1626908933
transform 1 0 7008 0 -1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_954
timestamp 1626908933
transform 1 0 7152 0 1 481
box -29 -23 29 23
use L1M1_PR  L1M1_PR_580
timestamp 1626908933
transform 1 0 7056 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_452
timestamp 1626908933
transform 1 0 7152 0 1 481
box -29 -23 29 23
use L1M1_PR  L1M1_PR_78
timestamp 1626908933
transform 1 0 7056 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_545
timestamp 1626908933
transform 1 0 7248 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_80
timestamp 1626908933
transform 1 0 7248 0 1 333
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_74
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_78
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_156
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_160
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_32
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_151
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_32
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_151
timestamp 1626908933
transform 1 0 7700 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_36
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_139
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_58
timestamp 1626908933
transform 1 0 7104 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_178
timestamp 1626908933
transform 1 0 7104 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_0
timestamp 1626908933
transform 1 0 7104 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_7
timestamp 1626908933
transform 1 0 7104 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_8
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_40
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 710 715
use M1M2_PR  M1M2_PR_662
timestamp 1626908933
transform 1 0 7920 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_197
timestamp 1626908933
transform 1 0 7920 0 1 407
box -32 -32 32 32
use L1M1_PR  L1M1_PR_246
timestamp 1626908933
transform 1 0 8688 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_476
timestamp 1626908933
transform 1 0 8592 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_748
timestamp 1626908933
transform 1 0 8688 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_978
timestamp 1626908933
transform 1 0 8592 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_251
timestamp 1626908933
transform 1 0 8304 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_434
timestamp 1626908933
transform 1 0 8496 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_716
timestamp 1626908933
transform 1 0 8304 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_899
timestamp 1626908933
transform 1 0 8496 0 1 407
box -32 -32 32 32
use L1M1_PR  L1M1_PR_303
timestamp 1626908933
transform 1 0 8400 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_805
timestamp 1626908933
transform 1 0 8400 0 1 555
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_0
timestamp 1626908933
transform 1 0 8256 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_2
timestamp 1626908933
transform 1 0 8256 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_7
timestamp 1626908933
transform -1 0 9024 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_39
timestamp 1626908933
transform -1 0 9024 0 1 0
box -38 -49 710 715
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_14
timestamp 1626908933
transform 1 0 8900 0 1 23
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_6
timestamp 1626908933
transform 1 0 8900 0 1 23
box -100 -26 100 26
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_14
timestamp 1626908933
transform 1 0 8900 0 1 16
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_6
timestamp 1626908933
transform 1 0 8900 0 1 16
box -100 -33 100 33
use L1M1_PR  L1M1_PR_953
timestamp 1626908933
transform 1 0 8976 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_451
timestamp 1626908933
transform 1 0 8976 0 1 111
box -29 -23 29 23
use L1M1_PR  L1M1_PR_576
timestamp 1626908933
transform 1 0 9072 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_74
timestamp 1626908933
transform 1 0 9072 0 1 555
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_154
timestamp 1626908933
transform 1 0 9024 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_147
timestamp 1626908933
transform 1 0 9024 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_41
timestamp 1626908933
transform 1 0 9024 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_34
timestamp 1626908933
transform 1 0 9024 0 1 0
box -38 -49 230 715
use M1M2_PR  M1M2_PR_73
timestamp 1626908933
transform 1 0 9552 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_538
timestamp 1626908933
transform 1 0 9552 0 1 555
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_30
timestamp 1626908933
transform 1 0 9216 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_133
timestamp 1626908933
transform 1 0 9216 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__and2b_2  sky130_fd_sc_hs__and2b_2_0
timestamp 1626908933
transform 1 0 9216 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__and2b_2  sky130_fd_sc_hs__and2b_2_1
timestamp 1626908933
transform 1 0 9216 0 -1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_155
timestamp 1626908933
transform 1 0 9888 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_42
timestamp 1626908933
transform 1 0 9888 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_159
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_77
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_38
timestamp 1626908933
transform 1 0 10080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_158
timestamp 1626908933
transform 1 0 10080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_39
timestamp 1626908933
transform 1 0 10464 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_152
timestamp 1626908933
transform 1 0 10464 0 1 0
box -38 -49 230 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_21
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_140
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_21
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_140
timestamp 1626908933
transform 1 0 10100 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_86
timestamp 1626908933
transform 1 0 10656 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_256
timestamp 1626908933
transform 1 0 10656 0 1 0
box -38 -49 134 715
use M1M2_PR  M1M2_PR_107
timestamp 1626908933
transform 1 0 10704 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_572
timestamp 1626908933
transform 1 0 10704 0 1 555
box -32 -32 32 32
use L1M1_PR  L1M1_PR_101
timestamp 1626908933
transform 1 0 10704 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_603
timestamp 1626908933
transform 1 0 10704 0 1 555
box -29 -23 29 23
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_2
timestamp 1626908933
transform 1 0 10752 0 1 0
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_3
timestamp 1626908933
transform -1 0 10560 0 -1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_8
timestamp 1626908933
transform 1 0 10752 0 1 0
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_9
timestamp 1626908933
transform -1 0 10560 0 -1 1332
box -38 -49 518 715
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_13
timestamp 1626908933
transform 1 0 11300 0 1 23
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_5
timestamp 1626908933
transform 1 0 11300 0 1 23
box -100 -26 100 26
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_13
timestamp 1626908933
transform 1 0 11300 0 1 16
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_5
timestamp 1626908933
transform 1 0 11300 0 1 16
box -100 -33 100 33
use L1M1_PR  L1M1_PR_970
timestamp 1626908933
transform 1 0 10992 0 1 259
box -29 -23 29 23
use L1M1_PR  L1M1_PR_468
timestamp 1626908933
transform 1 0 10992 0 1 259
box -29 -23 29 23
use L1M1_PR  L1M1_PR_779
timestamp 1626908933
transform 1 0 11184 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_277
timestamp 1626908933
transform 1 0 11184 0 1 555
box -29 -23 29 23
use M1M2_PR  M1M2_PR_692
timestamp 1626908933
transform 1 0 11472 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_227
timestamp 1626908933
transform 1 0 11472 0 1 555
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_145
timestamp 1626908933
transform 1 0 11232 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_25
timestamp 1626908933
transform 1 0 11232 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_82
timestamp 1626908933
transform 1 0 11616 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_252
timestamp 1626908933
transform 1 0 11616 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_17
timestamp 1626908933
transform 1 0 11712 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_120
timestamp 1626908933
transform 1 0 11712 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_72
timestamp 1626908933
transform -1 0 12480 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_35
timestamp 1626908933
transform -1 0 12480 0 -1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_73
timestamp 1626908933
transform 1 0 12480 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_76
timestamp 1626908933
transform 1 0 12480 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_155
timestamp 1626908933
transform 1 0 12480 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_158
timestamp 1626908933
transform 1 0 12480 0 1 0
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_10
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_129
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_10
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_129
timestamp 1626908933
transform 1 0 12500 0 1 666
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_14
timestamp 1626908933
transform 1 0 12576 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_15
timestamp 1626908933
transform 1 0 12576 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_134
timestamp 1626908933
transform 1 0 12576 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_135
timestamp 1626908933
transform 1 0 12576 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_112
timestamp 1626908933
transform 1 0 12960 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_111
timestamp 1626908933
transform 1 0 12960 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_9
timestamp 1626908933
transform 1 0 12960 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_8
timestamp 1626908933
transform 1 0 12960 0 -1 1332
box -38 -49 806 715
use M2M3_PR  M2M3_PR_48
timestamp 1626908933
transform 1 0 13776 0 1 281
box -33 -37 33 37
use M2M3_PR  M2M3_PR_6
timestamp 1626908933
transform 1 0 13776 0 1 281
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_258
timestamp 1626908933
transform 1 0 13920 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_257
timestamp 1626908933
transform 1 0 13920 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_88
timestamp 1626908933
transform 1 0 13920 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_87
timestamp 1626908933
transform 1 0 13920 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_156
timestamp 1626908933
transform 1 0 13728 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_153
timestamp 1626908933
transform 1 0 13728 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_43
timestamp 1626908933
transform 1 0 13728 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_40
timestamp 1626908933
transform 1 0 13728 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_72
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_154
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_44
timestamp 1626908933
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_157
timestamp 1626908933
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_89
timestamp 1626908933
transform 1 0 192 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_259
timestamp 1626908933
transform 1 0 192 0 1 1332
box -38 -49 134 715
use M2M3_PR  M2M3_PR_27
timestamp 1626908933
transform 1 0 240 0 1 1257
box -33 -37 33 37
use M2M3_PR  M2M3_PR_69
timestamp 1626908933
transform 1 0 240 0 1 1257
box -33 -37 33 37
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_91
timestamp 1626908933
transform 1 0 768 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_194
timestamp 1626908933
transform 1 0 768 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_118
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_238
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_418
timestamp 1626908933
transform 1 0 912 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_883
timestamp 1626908933
transform 1 0 912 0 1 1443
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_78
timestamp 1626908933
transform 1 0 1536 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_248
timestamp 1626908933
transform 1 0 1536 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_417
timestamp 1626908933
transform 1 0 1680 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_882
timestamp 1626908933
transform 1 0 1680 0 1 1221
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_118
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_237
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_118
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_237
timestamp 1626908933
transform 1 0 1700 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_102
timestamp 1626908933
transform 1 0 1632 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_222
timestamp 1626908933
transform 1 0 1632 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_260
timestamp 1626908933
transform 1 0 2112 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_247
timestamp 1626908933
transform 1 0 2016 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_90
timestamp 1626908933
transform 1 0 2112 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_77
timestamp 1626908933
transform 1 0 2016 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_881
timestamp 1626908933
transform 1 0 3312 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_554
timestamp 1626908933
transform 1 0 3888 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_416
timestamp 1626908933
transform 1 0 3312 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_89
timestamp 1626908933
transform 1 0 3888 0 1 777
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_46
timestamp 1626908933
transform 1 0 2208 0 1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_9
timestamp 1626908933
transform 1 0 2208 0 1 1332
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_588
timestamp 1626908933
transform 1 0 4272 0 1 777
box -29 -23 29 23
use L1M1_PR  L1M1_PR_86
timestamp 1626908933
transform 1 0 4272 0 1 777
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_227
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_108
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_227
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_108
timestamp 1626908933
transform 1 0 4100 0 1 1332
box -100 -49 100 49
use L1M1_PR  L1M1_PR_960
timestamp 1626908933
transform 1 0 4176 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_458
timestamp 1626908933
transform 1 0 4176 0 1 1443
box -29 -23 29 23
use M1M2_PR  M1M2_PR_910
timestamp 1626908933
transform 1 0 4368 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_445
timestamp 1626908933
transform 1 0 4368 0 1 1443
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_71
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_153
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_45
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_158
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 230 715
use M1M2_PR  M1M2_PR_244
timestamp 1626908933
transform 1 0 4560 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_709
timestamp 1626908933
transform 1 0 4560 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_0
timestamp 1626908933
transform 1 0 4128 0 1 1332
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_32
timestamp 1626908933
transform 1 0 4128 0 1 1332
box -38 -49 710 715
use L1M1_PR  L1M1_PR_798
timestamp 1626908933
transform 1 0 5616 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_296
timestamp 1626908933
transform 1 0 5616 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_548
timestamp 1626908933
transform 1 0 5136 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_83
timestamp 1626908933
transform 1 0 5136 0 1 1443
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_156
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_53
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_48
timestamp 1626908933
transform 1 0 5856 0 1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_11
timestamp 1626908933
transform 1 0 5856 0 1 1332
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_318
timestamp 1626908933
transform 1 0 6096 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_783
timestamp 1626908933
transform 1 0 6096 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_372
timestamp 1626908933
transform 1 0 6000 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_874
timestamp 1626908933
transform 1 0 6000 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_69
timestamp 1626908933
transform 1 0 6672 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_534
timestamp 1626908933
transform 1 0 6672 0 1 999
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_98
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_217
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_98
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_217
timestamp 1626908933
transform 1 0 6500 0 1 1332
box -100 -49 100 49
use M1M2_PR  M1M2_PR_79
timestamp 1626908933
transform 1 0 7248 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_408
timestamp 1626908933
transform 1 0 7056 0 1 1147
box -32 -32 32 32
use M1M2_PR  M1M2_PR_544
timestamp 1626908933
transform 1 0 7248 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_873
timestamp 1626908933
transform 1 0 7056 0 1 1147
box -32 -32 32 32
use L1M1_PR  L1M1_PR_80
timestamp 1626908933
transform 1 0 7440 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_582
timestamp 1626908933
transform 1 0 7440 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_46
timestamp 1626908933
transform 1 0 7776 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_159
timestamp 1626908933
transform 1 0 7776 0 1 1332
box -38 -49 230 715
use L1M1_PR  L1M1_PR_69
timestamp 1626908933
transform 1 0 7632 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_450
timestamp 1626908933
transform 1 0 7632 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_571
timestamp 1626908933
transform 1 0 7632 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_952
timestamp 1626908933
transform 1 0 7632 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_196
timestamp 1626908933
transform 1 0 7920 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_661
timestamp 1626908933
transform 1 0 7920 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_248
timestamp 1626908933
transform 1 0 7920 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_750
timestamp 1626908933
transform 1 0 7920 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_49
timestamp 1626908933
transform 1 0 7968 0 1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_12
timestamp 1626908933
transform 1 0 7968 0 1 1332
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_981
timestamp 1626908933
transform 1 0 8016 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_479
timestamp 1626908933
transform 1 0 8016 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_807
timestamp 1626908933
transform 1 0 8208 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_305
timestamp 1626908933
transform 1 0 8208 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_898
timestamp 1626908933
transform 1 0 8496 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_433
timestamp 1626908933
transform 1 0 8496 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_718
timestamp 1626908933
transform 1 0 8688 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_253
timestamp 1626908933
transform 1 0 8688 0 1 1221
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_207
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_88
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_207
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_88
timestamp 1626908933
transform 1 0 8900 0 1 1332
box -100 -49 100 49
use L1M1_PR  L1M1_PR_977
timestamp 1626908933
transform 1 0 8976 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_475
timestamp 1626908933
transform 1 0 8976 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_887
timestamp 1626908933
transform 1 0 9072 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_422
timestamp 1626908933
transform 1 0 9072 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_975
timestamp 1626908933
transform 1 0 9264 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_473
timestamp 1626908933
transform 1 0 9264 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_746
timestamp 1626908933
transform 1 0 9456 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_244
timestamp 1626908933
transform 1 0 9456 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_961
timestamp 1626908933
transform 1 0 9648 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_577
timestamp 1626908933
transform 1 0 9744 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_459
timestamp 1626908933
transform 1 0 9648 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_75
timestamp 1626908933
transform 1 0 9744 0 1 1443
box -29 -23 29 23
use M1M2_PR  M1M2_PR_541
timestamp 1626908933
transform 1 0 9744 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_540
timestamp 1626908933
transform 1 0 9744 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_76
timestamp 1626908933
transform 1 0 9744 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_75
timestamp 1626908933
transform 1 0 9744 0 1 1443
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_261
timestamp 1626908933
transform 1 0 9888 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_91
timestamp 1626908933
transform 1 0 9888 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_152
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_70
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_37
timestamp 1626908933
transform 1 0 10080 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_157
timestamp 1626908933
transform 1 0 10080 0 1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_279
timestamp 1626908933
transform 1 0 10224 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_470
timestamp 1626908933
transform 1 0 10320 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_781
timestamp 1626908933
transform 1 0 10224 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_972
timestamp 1626908933
transform 1 0 10320 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_602
timestamp 1626908933
transform 1 0 10704 0 1 777
box -29 -23 29 23
use L1M1_PR  L1M1_PR_100
timestamp 1626908933
transform 1 0 10704 0 1 777
box -29 -23 29 23
use M1M2_PR  M1M2_PR_571
timestamp 1626908933
transform 1 0 10704 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_106
timestamp 1626908933
transform 1 0 10704 0 1 777
box -32 -32 32 32
use L1M1_PR  L1M1_PR_605
timestamp 1626908933
transform 1 0 10512 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_103
timestamp 1626908933
transform 1 0 10512 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_694
timestamp 1626908933
transform 1 0 10608 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_574
timestamp 1626908933
transform 1 0 10704 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_229
timestamp 1626908933
transform 1 0 10608 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_109
timestamp 1626908933
transform 1 0 10704 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_604
timestamp 1626908933
transform 1 0 10608 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_102
timestamp 1626908933
transform 1 0 10608 0 1 1443
box -29 -23 29 23
use M1M2_PR  M1M2_PR_573
timestamp 1626908933
transform 1 0 10704 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_108
timestamp 1626908933
transform 1 0 10704 0 1 1443
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_197
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_78
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_197
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_78
timestamp 1626908933
transform 1 0 11300 0 1 1332
box -100 -49 100 49
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_71
timestamp 1626908933
transform -1 0 12384 0 1 1332
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_34
timestamp 1626908933
transform -1 0 12384 0 1 1332
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_224
timestamp 1626908933
transform 1 0 12144 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_225
timestamp 1626908933
transform 1 0 12144 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_689
timestamp 1626908933
transform 1 0 12144 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_690
timestamp 1626908933
transform 1 0 12144 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_275
timestamp 1626908933
transform 1 0 12048 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_777
timestamp 1626908933
transform 1 0 12048 0 1 1073
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_32
timestamp 1626908933
transform 1 0 12384 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_145
timestamp 1626908933
transform 1 0 12384 0 1 1332
box -38 -49 230 715
use M1M2_PR  M1M2_PR_295
timestamp 1626908933
transform 1 0 12336 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_760
timestamp 1626908933
transform 1 0 12336 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_353
timestamp 1626908933
transform 1 0 12432 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_855
timestamp 1626908933
transform 1 0 12432 0 1 999
box -29 -23 29 23
use M1M2_PR  M1M2_PR_398
timestamp 1626908933
transform 1 0 12528 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_863
timestamp 1626908933
transform 1 0 12528 0 1 777
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_7
timestamp 1626908933
transform -1 0 13536 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_1
timestamp 1626908933
transform -1 0 13536 0 1 1332
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_246
timestamp 1626908933
transform 1 0 12576 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_76
timestamp 1626908933
transform 1 0 12576 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_133
timestamp 1626908933
transform 1 0 12672 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_13
timestamp 1626908933
transform 1 0 12672 0 1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_274
timestamp 1626908933
transform 1 0 13200 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_776
timestamp 1626908933
transform 1 0 13200 0 1 1443
box -29 -23 29 23
use M2M3_PR  M2M3_PR_5
timestamp 1626908933
transform 1 0 13488 0 1 891
box -33 -37 33 37
use M2M3_PR  M2M3_PR_47
timestamp 1626908933
transform 1 0 13488 0 1 891
box -33 -37 33 37
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_69
timestamp 1626908933
transform 1 0 13632 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_151
timestamp 1626908933
transform 1 0 13632 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_92
timestamp 1626908933
transform 1 0 13536 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_262
timestamp 1626908933
transform 1 0 13536 0 1 1332
box -38 -49 134 715
use prbs_generator_syn_VIA8  prbs_generator_syn_VIA8_0
timestamp 1626908933
transform 1 0 13700 0 1 1317
box -100 -34 100 34
use prbs_generator_syn_VIA8  prbs_generator_syn_VIA8_1
timestamp 1626908933
transform 1 0 13700 0 1 1317
box -100 -34 100 34
use prbs_generator_syn_VIA9  prbs_generator_syn_VIA9_0
timestamp 1626908933
transform 1 0 13700 0 1 1317
box -100 -34 100 34
use prbs_generator_syn_VIA9  prbs_generator_syn_VIA9_1
timestamp 1626908933
transform 1 0 13700 0 1 1317
box -100 -34 100 34
use M2M3_PR  M2M3_PR_49
timestamp 1626908933
transform 1 0 13776 0 1 1501
box -33 -37 33 37
use M2M3_PR  M2M3_PR_7
timestamp 1626908933
transform 1 0 13776 0 1 1501
box -33 -37 33 37
use M1M2_PR  M1M2_PR_862
timestamp 1626908933
transform 1 0 13968 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_397
timestamp 1626908933
transform 1 0 13968 0 1 777
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_263
timestamp 1626908933
transform 1 0 13920 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_93
timestamp 1626908933
transform 1 0 13920 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_160
timestamp 1626908933
transform 1 0 13728 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_47
timestamp 1626908933
transform 1 0 13728 0 1 1332
box -38 -49 230 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_183
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_64
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_183
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_64
timestamp 1626908933
transform 1 0 500 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_245
timestamp 1626908933
transform 1 0 0 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_75
timestamp 1626908933
transform 1 0 0 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_204
timestamp 1626908933
transform 1 0 96 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_101
timestamp 1626908933
transform 1 0 96 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_244
timestamp 1626908933
transform 1 0 1248 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_74
timestamp 1626908933
transform 1 0 1248 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_229
timestamp 1626908933
transform 1 0 864 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_109
timestamp 1626908933
transform 1 0 864 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_184
timestamp 1626908933
transform 1 0 1344 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_81
timestamp 1626908933
transform 1 0 1344 0 -1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_95
timestamp 1626908933
transform 1 0 2256 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_560
timestamp 1626908933
transform 1 0 2256 0 1 1887
box -32 -32 32 32
use L1M1_PR  L1M1_PR_388
timestamp 1626908933
transform 1 0 2256 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_890
timestamp 1626908933
transform 1 0 2256 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_150
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_68
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_797
timestamp 1626908933
transform 1 0 2640 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_295
timestamp 1626908933
transform 1 0 2640 0 1 1591
box -29 -23 29 23
use M1M2_PR  M1M2_PR_707
timestamp 1626908933
transform 1 0 2640 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_242
timestamp 1626908933
transform 1 0 2640 0 1 1591
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_172
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_53
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_172
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_53
timestamp 1626908933
transform 1 0 2900 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_70
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_173
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_94
timestamp 1626908933
transform 1 0 2112 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_214
timestamp 1626908933
transform 1 0 2112 0 -1 2664
box -38 -49 422 715
use M1M2_PR  M1M2_PR_797
timestamp 1626908933
transform 1 0 3120 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_332
timestamp 1626908933
transform 1 0 3120 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_144
timestamp 1626908933
transform 1 0 3360 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_31
timestamp 1626908933
transform 1 0 3360 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_164
timestamp 1626908933
transform 1 0 3552 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_61
timestamp 1626908933
transform 1 0 3552 0 -1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_591
timestamp 1626908933
transform 1 0 3792 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_89
timestamp 1626908933
transform 1 0 3792 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_96
timestamp 1626908933
transform 1 0 4272 0 1 1675
box -29 -23 29 23
use L1M1_PR  L1M1_PR_598
timestamp 1626908933
transform 1 0 4272 0 1 1675
box -29 -23 29 23
use M1M2_PR  M1M2_PR_100
timestamp 1626908933
transform 1 0 4464 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_205
timestamp 1626908933
transform 1 0 4464 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_565
timestamp 1626908933
transform 1 0 4464 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_670
timestamp 1626908933
transform 1 0 4464 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_256
timestamp 1626908933
transform 1 0 4464 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_758
timestamp 1626908933
transform 1 0 4464 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_486
timestamp 1626908933
transform 1 0 4578 0 1 1619
box -29 -23 29 23
use L1M1_PR  L1M1_PR_988
timestamp 1626908933
transform 1 0 4578 0 1 1619
box -29 -23 29 23
use L1M1_PR  L1M1_PR_373
timestamp 1626908933
transform 1 0 5904 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_875
timestamp 1626908933
transform 1 0 5904 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_87
timestamp 1626908933
transform 1 0 4272 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_552
timestamp 1626908933
transform 1 0 4272 0 1 2109
box -32 -32 32 32
use L1M1_PR  L1M1_PR_83
timestamp 1626908933
transform 1 0 4464 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_585
timestamp 1626908933
transform 1 0 4464 0 1 2109
box -29 -23 29 23
use M1M2_PR  M1M2_PR_202
timestamp 1626908933
transform 1 0 4752 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_667
timestamp 1626908933
transform 1 0 4752 0 1 2257
box -32 -32 32 32
use L1M1_PR  L1M1_PR_289
timestamp 1626908933
transform 1 0 4752 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_791
timestamp 1626908933
transform 1 0 4752 0 1 1887
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_42
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_161
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_42
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_161
timestamp 1626908933
transform 1 0 5300 0 1 1998
box -100 -49 100 49
use M1M2_PR  M1M2_PR_86
timestamp 1626908933
transform 1 0 5616 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_551
timestamp 1626908933
transform 1 0 5616 0 1 2109
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_47
timestamp 1626908933
transform -1 0 6240 0 -1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_10
timestamp 1626908933
transform -1 0 6240 0 -1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_73
timestamp 1626908933
transform 1 0 6240 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_243
timestamp 1626908933
transform 1 0 6240 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_248
timestamp 1626908933
transform 1 0 6288 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_317
timestamp 1626908933
transform 1 0 6096 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_713
timestamp 1626908933
transform 1 0 6288 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_782
timestamp 1626908933
transform 1 0 6096 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_301
timestamp 1626908933
transform 1 0 6288 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_803
timestamp 1626908933
transform 1 0 6288 0 1 1591
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_63
timestamp 1626908933
transform 1 0 6336 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_183
timestamp 1626908933
transform 1 0 6336 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_9
timestamp 1626908933
transform -1 0 7392 0 -1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_41
timestamp 1626908933
transform -1 0 7392 0 -1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_264
timestamp 1626908933
transform 1 0 7392 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_94
timestamp 1626908933
transform 1 0 7392 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_149
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_67
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_72
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_242
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_31
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_150
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_31
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_150
timestamp 1626908933
transform 1 0 7700 0 1 1998
box -100 -49 100 49
use M1M2_PR  M1M2_PR_313
timestamp 1626908933
transform 1 0 7920 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_778
timestamp 1626908933
transform 1 0 7920 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_54
timestamp 1626908933
transform 1 0 7680 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_174
timestamp 1626908933
transform 1 0 7680 0 -1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_366
timestamp 1626908933
transform 1 0 8016 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_868
timestamp 1626908933
transform 1 0 8016 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_250
timestamp 1626908933
transform 1 0 8304 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_715
timestamp 1626908933
transform 1 0 8304 0 1 1591
box -32 -32 32 32
use L1M1_PR  L1M1_PR_302
timestamp 1626908933
transform 1 0 8400 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_804
timestamp 1626908933
transform 1 0 8400 0 1 1591
box -29 -23 29 23
use M1M2_PR  M1M2_PR_239
timestamp 1626908933
transform 1 0 8304 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_704
timestamp 1626908933
transform 1 0 8304 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_77
timestamp 1626908933
transform 1 0 8880 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_542
timestamp 1626908933
transform 1 0 8880 0 1 1813
box -32 -32 32 32
use M1M2_PR  M1M2_PR_421
timestamp 1626908933
transform 1 0 9072 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_886
timestamp 1626908933
transform 1 0 9072 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_72
timestamp 1626908933
transform 1 0 9552 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_537
timestamp 1626908933
transform 1 0 9552 0 1 2109
box -32 -32 32 32
use L1M1_PR  L1M1_PR_72
timestamp 1626908933
transform 1 0 9648 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_76
timestamp 1626908933
transform 1 0 9552 0 1 1813
box -29 -23 29 23
use L1M1_PR  L1M1_PR_574
timestamp 1626908933
transform 1 0 9648 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_578
timestamp 1626908933
transform 1 0 9552 0 1 1813
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_71
timestamp 1626908933
transform 1 0 9984 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_241
timestamp 1626908933
transform 1 0 9984 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_82
timestamp 1626908933
transform 1 0 9936 0 1 1517
box -32 -32 32 32
use M1M2_PR  M1M2_PR_547
timestamp 1626908933
transform 1 0 9936 0 1 1517
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_50
timestamp 1626908933
transform 1 0 8064 0 -1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_13
timestamp 1626908933
transform 1 0 8064 0 -1 2664
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_139
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_20
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_139
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_20
timestamp 1626908933
transform 1 0 10100 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_240
timestamp 1626908933
transform 1 0 10464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_70
timestamp 1626908933
transform 1 0 10464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_156
timestamp 1626908933
transform 1 0 10080 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_36
timestamp 1626908933
transform 1 0 10080 0 -1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_778
timestamp 1626908933
transform 1 0 11952 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_276
timestamp 1626908933
transform 1 0 11952 0 1 1591
box -29 -23 29 23
use M1M2_PR  M1M2_PR_761
timestamp 1626908933
transform 1 0 11760 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_691
timestamp 1626908933
transform 1 0 11472 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_296
timestamp 1626908933
transform 1 0 11760 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_226
timestamp 1626908933
transform 1 0 11472 0 1 1591
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_70
timestamp 1626908933
transform 1 0 10560 0 -1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_33
timestamp 1626908933
transform 1 0 10560 0 -1 2664
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_294
timestamp 1626908933
transform 1 0 12336 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_759
timestamp 1626908933
transform 1 0 12336 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_354
timestamp 1626908933
transform 1 0 12336 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_856
timestamp 1626908933
transform 1 0 12336 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_66
timestamp 1626908933
transform 1 0 12480 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_148
timestamp 1626908933
transform 1 0 12480 0 -1 2664
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_9
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_128
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_9
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_128
timestamp 1626908933
transform 1 0 12500 0 1 1998
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_12
timestamp 1626908933
transform 1 0 12576 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_132
timestamp 1626908933
transform 1 0 12576 0 -1 2664
box -38 -49 422 715
use L1M1_PR  L1M1_PR_963
timestamp 1626908933
transform 1 0 13296 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_896
timestamp 1626908933
transform 1 0 13584 0 1 1517
box -29 -23 29 23
use L1M1_PR  L1M1_PR_461
timestamp 1626908933
transform 1 0 13296 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_394
timestamp 1626908933
transform 1 0 13584 0 1 1517
box -29 -23 29 23
use M1M2_PR  M1M2_PR_890
timestamp 1626908933
transform 1 0 12912 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_425
timestamp 1626908933
transform 1 0 12912 0 1 1591
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_110
timestamp 1626908933
transform 1 0 12960 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_7
timestamp 1626908933
transform 1 0 12960 0 -1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_884
timestamp 1626908933
transform 1 0 13680 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_803
timestamp 1626908933
transform 1 0 13776 0 1 1517
box -32 -32 32 32
use M1M2_PR  M1M2_PR_419
timestamp 1626908933
transform 1 0 13680 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_338
timestamp 1626908933
transform 1 0 13776 0 1 1517
box -32 -32 32 32
use M2M3_PR  M2M3_PR_82
timestamp 1626908933
transform 1 0 13680 0 1 2111
box -33 -37 33 37
use M2M3_PR  M2M3_PR_40
timestamp 1626908933
transform 1 0 13680 0 1 2111
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_265
timestamp 1626908933
transform 1 0 13920 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_95
timestamp 1626908933
transform 1 0 13920 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_161
timestamp 1626908933
transform 1 0 13728 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_48
timestamp 1626908933
transform 1 0 13728 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_65
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_147
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_49
timestamp 1626908933
transform 1 0 0 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_162
timestamp 1626908933
transform 1 0 0 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_96
timestamp 1626908933
transform 1 0 192 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_266
timestamp 1626908933
transform 1 0 192 0 1 2664
box -38 -49 134 715
use M2M3_PR  M2M3_PR_28
timestamp 1626908933
transform 1 0 240 0 1 2355
box -33 -37 33 37
use M2M3_PR  M2M3_PR_70
timestamp 1626908933
transform 1 0 240 0 1 2355
box -33 -37 33 37
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_90
timestamp 1626908933
transform 1 0 768 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_193
timestamp 1626908933
transform 1 0 768 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_117
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_237
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 422 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_236
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_117
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_236
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_117
timestamp 1626908933
transform 1 0 1700 0 1 2664
box -100 -49 100 49
use M1M2_PR  M1M2_PR_926
timestamp 1626908933
transform 1 0 1488 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_461
timestamp 1626908933
transform 1 0 1488 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_267
timestamp 1626908933
transform 1 0 1536 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_97
timestamp 1626908933
transform 1 0 1536 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_795
timestamp 1626908933
transform 1 0 1680 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_293
timestamp 1626908933
transform 1 0 1680 0 1 2923
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_2
timestamp 1626908933
transform -1 0 2304 0 1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_34
timestamp 1626908933
transform -1 0 2304 0 1 2664
box -38 -49 710 715
use L1M1_PR  L1M1_PR_996
timestamp 1626908933
transform 1 0 1872 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_764
timestamp 1626908933
transform 1 0 1968 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_494
timestamp 1626908933
transform 1 0 1872 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_262
timestamp 1626908933
transform 1 0 1968 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_674
timestamp 1626908933
transform 1 0 1968 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_209
timestamp 1626908933
transform 1 0 1968 0 1 2997
box -32 -32 32 32
use L1M1_PR  L1M1_PR_958
timestamp 1626908933
transform 1 0 2256 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_592
timestamp 1626908933
transform 1 0 2256 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_456
timestamp 1626908933
transform 1 0 2256 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_90
timestamp 1626908933
transform 1 0 2256 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_879
timestamp 1626908933
transform 1 0 2448 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_559
timestamp 1626908933
transform 1 0 2256 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_414
timestamp 1626908933
transform 1 0 2448 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_94
timestamp 1626908933
transform 1 0 2256 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_213
timestamp 1626908933
transform 1 0 2304 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_93
timestamp 1626908933
transform 1 0 2304 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_50
timestamp 1626908933
transform 1 0 2688 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_163
timestamp 1626908933
transform 1 0 2688 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_98
timestamp 1626908933
transform 1 0 2880 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_268
timestamp 1626908933
transform 1 0 2880 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_886
timestamp 1626908933
transform 1 0 3024 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_794
timestamp 1626908933
transform 1 0 3408 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_384
timestamp 1626908933
transform 1 0 3024 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_292
timestamp 1626908933
transform 1 0 3408 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_796
timestamp 1626908933
transform 1 0 3120 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_794
timestamp 1626908933
transform 1 0 3504 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_331
timestamp 1626908933
transform 1 0 3120 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_329
timestamp 1626908933
transform 1 0 3504 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_45
timestamp 1626908933
transform 1 0 2976 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_8
timestamp 1626908933
transform 1 0 2976 0 1 2664
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_226
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_107
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_226
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_107
timestamp 1626908933
transform 1 0 4100 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_269
timestamp 1626908933
transform 1 0 4896 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_99
timestamp 1626908933
transform 1 0 4896 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_146
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_64
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_801
timestamp 1626908933
transform 1 0 5808 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_299
timestamp 1626908933
transform 1 0 5808 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_711
timestamp 1626908933
transform 1 0 5904 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_246
timestamp 1626908933
transform 1 0 5904 0 1 2331
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_270
timestamp 1626908933
transform 1 0 5280 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_100
timestamp 1626908933
transform 1 0 5280 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_164
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_51
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_51
timestamp 1626908933
transform -1 0 7296 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_14
timestamp 1626908933
transform -1 0 7296 0 1 2664
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_316
timestamp 1626908933
transform 1 0 6096 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_781
timestamp 1626908933
transform 1 0 6096 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_371
timestamp 1626908933
transform 1 0 6192 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_873
timestamp 1626908933
transform 1 0 6192 0 1 2331
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_97
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_216
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_97
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_216
timestamp 1626908933
transform 1 0 6500 0 1 2664
box -100 -49 100 49
use M1M2_PR  M1M2_PR_255
timestamp 1626908933
transform 1 0 6672 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_720
timestamp 1626908933
transform 1 0 6672 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_307
timestamp 1626908933
transform 1 0 6768 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_809
timestamp 1626908933
transform 1 0 6768 0 1 2553
box -29 -23 29 23
use M1M2_PR  M1M2_PR_254
timestamp 1626908933
transform 1 0 6672 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_719
timestamp 1626908933
transform 1 0 6672 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_983
timestamp 1626908933
transform 1 0 6960 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_481
timestamp 1626908933
transform 1 0 6960 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_905
timestamp 1626908933
transform 1 0 6960 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_440
timestamp 1626908933
transform 1 0 6960 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_752
timestamp 1626908933
transform 1 0 7056 0 1 2321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_250
timestamp 1626908933
transform 1 0 7056 0 1 2321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_569
timestamp 1626908933
transform 1 0 7248 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_67
timestamp 1626908933
transform 1 0 7248 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_533
timestamp 1626908933
transform 1 0 7248 0 1 2479
box -32 -32 32 32
use M1M2_PR  M1M2_PR_68
timestamp 1626908933
transform 1 0 7248 0 1 2479
box -32 -32 32 32
use L1M1_PR  L1M1_PR_808
timestamp 1626908933
transform 1 0 6864 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_306
timestamp 1626908933
transform 1 0 6864 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_904
timestamp 1626908933
transform 1 0 7056 0 1 2849
box -32 -32 32 32
use M1M2_PR  M1M2_PR_439
timestamp 1626908933
transform 1 0 7056 0 1 2849
box -32 -32 32 32
use L1M1_PR  L1M1_PR_872
timestamp 1626908933
transform 1 0 7248 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_370
timestamp 1626908933
transform 1 0 7248 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_69
timestamp 1626908933
transform 1 0 7296 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_239
timestamp 1626908933
transform 1 0 7296 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_407
timestamp 1626908933
transform 1 0 7536 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_438
timestamp 1626908933
transform 1 0 7440 0 1 2849
box -32 -32 32 32
use M1M2_PR  M1M2_PR_872
timestamp 1626908933
transform 1 0 7536 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_903
timestamp 1626908933
transform 1 0 7440 0 1 2849
box -32 -32 32 32
use L1M1_PR  L1M1_PR_449
timestamp 1626908933
transform 1 0 7344 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_951
timestamp 1626908933
transform 1 0 7344 0 1 2553
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_38
timestamp 1626908933
transform 1 0 7392 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_141
timestamp 1626908933
transform 1 0 7392 0 1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_777
timestamp 1626908933
transform 1 0 7920 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_776
timestamp 1626908933
transform 1 0 7920 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_312
timestamp 1626908933
transform 1 0 7920 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_311
timestamp 1626908933
transform 1 0 7920 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_252
timestamp 1626908933
transform 1 0 8688 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_717
timestamp 1626908933
transform 1 0 8688 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_304
timestamp 1626908933
transform 1 0 8496 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_365
timestamp 1626908933
transform 1 0 8112 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_806
timestamp 1626908933
transform 1 0 8496 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_867
timestamp 1626908933
transform 1 0 8112 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_432
timestamp 1626908933
transform 1 0 8496 0 1 2849
box -32 -32 32 32
use M1M2_PR  M1M2_PR_897
timestamp 1626908933
transform 1 0 8496 0 1 2849
box -32 -32 32 32
use L1M1_PR  L1M1_PR_460
timestamp 1626908933
transform 1 0 8592 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_477
timestamp 1626908933
transform 1 0 8400 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_962
timestamp 1626908933
transform 1 0 8592 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_979
timestamp 1626908933
transform 1 0 8400 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_32
timestamp 1626908933
transform 1 0 8640 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_135
timestamp 1626908933
transform 1 0 8640 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_0
timestamp 1626908933
transform -1 0 8640 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_1
timestamp 1626908933
transform -1 0 8640 0 1 2664
box -38 -49 518 715
use M1M2_PR  M1M2_PR_420
timestamp 1626908933
transform 1 0 9072 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_885
timestamp 1626908933
transform 1 0 9072 0 1 2923
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_87
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_206
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_87
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_206
timestamp 1626908933
transform 1 0 8900 0 1 2664
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_30
timestamp 1626908933
transform 1 0 9408 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_143
timestamp 1626908933
transform 1 0 9408 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_42
timestamp 1626908933
transform 1 0 9600 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_162
timestamp 1626908933
transform 1 0 9600 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_145
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_63
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_305
timestamp 1626908933
transform 1 0 10320 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_770
timestamp 1626908933
transform 1 0 10320 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_360
timestamp 1626908933
transform 1 0 10608 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_862
timestamp 1626908933
transform 1 0 10608 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_231
timestamp 1626908933
transform 1 0 11088 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_696
timestamp 1626908933
transform 1 0 11088 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_281
timestamp 1626908933
transform 1 0 10992 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_783
timestamp 1626908933
transform 1 0 10992 0 1 2331
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_77
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_196
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_77
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_196
timestamp 1626908933
transform 1 0 11300 0 1 2664
box -100 -49 100 49
use L1M1_PR  L1M1_PR_361
timestamp 1626908933
transform 1 0 10128 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_863
timestamp 1626908933
transform 1 0 10128 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_304
timestamp 1626908933
transform 1 0 10320 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_769
timestamp 1626908933
transform 1 0 10320 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_228
timestamp 1626908933
transform 1 0 10608 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_693
timestamp 1626908933
transform 1 0 10608 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_278
timestamp 1626908933
transform 1 0 10512 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_780
timestamp 1626908933
transform 1 0 10512 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_230
timestamp 1626908933
transform 1 0 11088 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_695
timestamp 1626908933
transform 1 0 11088 0 1 2775
box -32 -32 32 32
use L1M1_PR  L1M1_PR_106
timestamp 1626908933
transform 1 0 11856 0 1 2849
box -29 -23 29 23
use L1M1_PR  L1M1_PR_608
timestamp 1626908933
transform 1 0 11856 0 1 2849
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_69
timestamp 1626908933
transform 1 0 10080 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_32
timestamp 1626908933
transform 1 0 10080 0 1 2664
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_111
timestamp 1626908933
transform 1 0 12240 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_576
timestamp 1626908933
transform 1 0 12240 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_108
timestamp 1626908933
transform 1 0 12144 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_610
timestamp 1626908933
transform 1 0 12144 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_607
timestamp 1626908933
transform 1 0 12048 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_105
timestamp 1626908933
transform 1 0 12048 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_609
timestamp 1626908933
transform 1 0 12240 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_107
timestamp 1626908933
transform 1 0 12240 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_575
timestamp 1626908933
transform 1 0 12240 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_110
timestamp 1626908933
transform 1 0 12240 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_606
timestamp 1626908933
transform 1 0 12528 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_104
timestamp 1626908933
transform 1 0 12528 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_966
timestamp 1626908933
transform 1 0 12720 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_464
timestamp 1626908933
transform 1 0 12720 0 1 2923
box -29 -23 29 23
use M1M2_PR  M1M2_PR_566
timestamp 1626908933
transform 1 0 12144 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_101
timestamp 1626908933
transform 1 0 12144 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_0
timestamp 1626908933
transform 1 0 12000 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_4
timestamp 1626908933
transform 1 0 12480 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_6
timestamp 1626908933
transform 1 0 12000 0 1 2664
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_10
timestamp 1626908933
transform 1 0 12480 0 1 2664
box -38 -49 518 715
use L1M1_PR  L1M1_PR_782
timestamp 1626908933
transform 1 0 12816 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_280
timestamp 1626908933
transform 1 0 12816 0 1 2775
box -29 -23 29 23
use M2M3_PR  M2M3_PR_83
timestamp 1626908933
transform 1 0 12912 0 1 2721
box -33 -37 33 37
use M2M3_PR  M2M3_PR_41
timestamp 1626908933
transform 1 0 12912 0 1 2721
box -33 -37 33 37
use M1M2_PR  M1M2_PR_891
timestamp 1626908933
transform 1 0 12816 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_426
timestamp 1626908933
transform 1 0 12816 0 1 2923
box -32 -32 32 32
use L1M1_PR  L1M1_PR_895
timestamp 1626908933
transform 1 0 13392 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_599
timestamp 1626908933
transform 1 0 13296 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_393
timestamp 1626908933
transform 1 0 13392 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_97
timestamp 1626908933
transform 1 0 13296 0 1 2997
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_33
timestamp 1626908933
transform -1 0 13632 0 1 2664
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_67
timestamp 1626908933
transform -1 0 13632 0 1 2664
box -38 -49 710 715
use M1M2_PR  M1M2_PR_802
timestamp 1626908933
transform 1 0 13872 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_337
timestamp 1626908933
transform 1 0 13872 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_271
timestamp 1626908933
transform 1 0 13920 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_101
timestamp 1626908933
transform 1 0 13920 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_165
timestamp 1626908933
transform 1 0 13728 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_52
timestamp 1626908933
transform 1 0 13728 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_144
timestamp 1626908933
transform 1 0 13632 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_62
timestamp 1626908933
transform 1 0 13632 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_68
timestamp 1626908933
transform 1 0 0 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_238
timestamp 1626908933
transform 1 0 0 0 -1 3996
box -38 -49 134 715
use M2M3_PR  M2M3_PR_29
timestamp 1626908933
transform 1 0 240 0 1 3453
box -33 -37 33 37
use M2M3_PR  M2M3_PR_71
timestamp 1626908933
transform 1 0 240 0 1 3453
box -33 -37 33 37
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_63
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_182
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_63
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_182
timestamp 1626908933
transform 1 0 500 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_100
timestamp 1626908933
transform 1 0 96 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_203
timestamp 1626908933
transform 1 0 96 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_67
timestamp 1626908933
transform 1 0 864 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_102
timestamp 1626908933
transform 1 0 960 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_237
timestamp 1626908933
transform 1 0 864 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_272
timestamp 1626908933
transform 1 0 960 0 -1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_219
timestamp 1626908933
transform 1 0 1104 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_684
timestamp 1626908933
transform 1 0 1104 0 1 3737
box -32 -32 32 32
use L1M1_PR  L1M1_PR_4
timestamp 1626908933
transform 1 0 1200 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_506
timestamp 1626908933
transform 1 0 1200 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_5
timestamp 1626908933
transform 1 0 1296 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_460
timestamp 1626908933
transform 1 0 1488 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_470
timestamp 1626908933
transform 1 0 1296 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_925
timestamp 1626908933
transform 1 0 1488 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_268
timestamp 1626908933
transform 1 0 1392 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_499
timestamp 1626908933
transform 1 0 1488 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_770
timestamp 1626908933
transform 1 0 1392 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1001
timestamp 1626908933
transform 1 0 1488 0 1 3663
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_30
timestamp 1626908933
transform 1 0 1056 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_62
timestamp 1626908933
transform 1 0 1056 0 -1 3996
box -38 -49 710 715
use M1M2_PR  M1M2_PR_673
timestamp 1626908933
transform 1 0 1968 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_208
timestamp 1626908933
transform 1 0 1968 0 1 3589
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_179
timestamp 1626908933
transform 1 0 1728 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_76
timestamp 1626908933
transform 1 0 1728 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_61
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_143
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_387
timestamp 1626908933
transform 1 0 2640 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_889
timestamp 1626908933
transform 1 0 2640 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_241
timestamp 1626908933
transform 1 0 2928 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_706
timestamp 1626908933
transform 1 0 2928 0 1 3737
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_52
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_171
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_52
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_171
timestamp 1626908933
transform 1 0 2900 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_793
timestamp 1626908933
transform 1 0 3024 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_291
timestamp 1626908933
transform 1 0 3024 0 1 3737
box -29 -23 29 23
use M1M2_PR  M1M2_PR_795
timestamp 1626908933
transform 1 0 3408 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_563
timestamp 1626908933
transform 1 0 3696 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_562
timestamp 1626908933
transform 1 0 3696 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_330
timestamp 1626908933
transform 1 0 3408 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_98
timestamp 1626908933
transform 1 0 3696 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_97
timestamp 1626908933
transform 1 0 3696 0 1 3737
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_44
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_7
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_597
timestamp 1626908933
transform 1 0 4368 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_594
timestamp 1626908933
transform 1 0 4560 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_95
timestamp 1626908933
transform 1 0 4368 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_92
timestamp 1626908933
transform 1 0 4560 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_564
timestamp 1626908933
transform 1 0 4464 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_99
timestamp 1626908933
transform 1 0 4464 0 1 3441
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_158
timestamp 1626908933
transform 1 0 4512 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_55
timestamp 1626908933
transform 1 0 4512 0 -1 3996
box -38 -49 806 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_41
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_160
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_41
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_160
timestamp 1626908933
transform 1 0 5300 0 1 3330
box -100 -49 100 49
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_1
timestamp 1626908933
transform 1 0 5280 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_0
timestamp 1626908933
transform 1 0 5280 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_66
timestamp 1626908933
transform 1 0 5568 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_236
timestamp 1626908933
transform 1 0 5568 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_66
timestamp 1626908933
transform 1 0 5664 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_186
timestamp 1626908933
transform 1 0 5664 0 -1 3996
box -38 -49 422 715
use L1M1_PR  L1M1_PR_573
timestamp 1626908933
transform 1 0 5712 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_71
timestamp 1626908933
transform 1 0 5712 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_596
timestamp 1626908933
transform 1 0 6192 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_94
timestamp 1626908933
transform 1 0 6192 0 1 3441
box -29 -23 29 23
use M1M2_PR  M1M2_PR_536
timestamp 1626908933
transform 1 0 6000 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_71
timestamp 1626908933
transform 1 0 6000 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_273
timestamp 1626908933
transform 1 0 6144 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_235
timestamp 1626908933
transform 1 0 6048 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_103
timestamp 1626908933
transform 1 0 6144 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_65
timestamp 1626908933
transform 1 0 6048 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_31
timestamp 1626908933
transform 1 0 6240 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_2
timestamp 1626908933
transform 1 0 6240 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_29
timestamp 1626908933
transform 1 0 6528 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_142
timestamp 1626908933
transform 1 0 6528 0 -1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_93
timestamp 1626908933
transform 1 0 6672 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_558
timestamp 1626908933
transform 1 0 6672 0 1 3071
box -32 -32 32 32
use L1M1_PR  L1M1_PR_425
timestamp 1626908933
transform 1 0 6576 0 1 3441
box -29 -23 29 23
use L1M1_PR  L1M1_PR_927
timestamp 1626908933
transform 1 0 6576 0 1 3441
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_43
timestamp 1626908933
transform 1 0 6720 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_146
timestamp 1626908933
transform 1 0 6720 0 -1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_201
timestamp 1626908933
transform 1 0 7152 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_235
timestamp 1626908933
transform 1 0 7056 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_666
timestamp 1626908933
transform 1 0 7152 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_700
timestamp 1626908933
transform 1 0 7056 0 1 3219
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_60
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_142
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_437
timestamp 1626908933
transform 1 0 7440 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_902
timestamp 1626908933
transform 1 0 7440 0 1 3589
box -32 -32 32 32
use L1M1_PR  L1M1_PR_369
timestamp 1626908933
transform 1 0 7632 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_871
timestamp 1626908933
transform 1 0 7632 0 1 3663
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_30
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_149
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_30
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_149
timestamp 1626908933
transform 1 0 7700 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_310
timestamp 1626908933
transform 1 0 7920 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_775
timestamp 1626908933
transform 1 0 7920 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_43
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_6
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_790
timestamp 1626908933
transform 1 0 8016 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_786
timestamp 1626908933
transform 1 0 8208 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_288
timestamp 1626908933
transform 1 0 8016 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_284
timestamp 1626908933
transform 1 0 8208 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_703
timestamp 1626908933
transform 1 0 8304 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_238
timestamp 1626908933
transform 1 0 8304 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_601
timestamp 1626908933
transform 1 0 9168 0 1 3515
box -29 -23 29 23
use L1M1_PR  L1M1_PR_99
timestamp 1626908933
transform 1 0 9168 0 1 3515
box -29 -23 29 23
use M1M2_PR  M1M2_PR_570
timestamp 1626908933
transform 1 0 9168 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_569
timestamp 1626908933
transform 1 0 9168 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_105
timestamp 1626908933
transform 1 0 9168 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_104
timestamp 1626908933
transform 1 0 9168 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_193
timestamp 1626908933
transform 1 0 9840 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_195
timestamp 1626908933
transform 1 0 9648 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_658
timestamp 1626908933
transform 1 0 9840 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_660
timestamp 1626908933
transform 1 0 9648 0 1 3589
box -32 -32 32 32
use L1M1_PR  L1M1_PR_243
timestamp 1626908933
transform 1 0 9840 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_472
timestamp 1626908933
transform 1 0 9744 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_745
timestamp 1626908933
transform 1 0 9840 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_974
timestamp 1626908933
transform 1 0 9744 0 1 3663
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_11
timestamp 1626908933
transform -1 0 10176 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_43
timestamp 1626908933
transform -1 0 10176 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_104
timestamp 1626908933
transform 1 0 10176 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_274
timestamp 1626908933
transform 1 0 10176 0 -1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_430
timestamp 1626908933
transform 1 0 10128 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_895
timestamp 1626908933
transform 1 0 10128 0 1 3515
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_19
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_138
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_19
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_138
timestamp 1626908933
transform 1 0 10100 0 1 3330
box -100 -49 100 49
use M1M2_PR  M1M2_PR_893
timestamp 1626908933
transform 1 0 10704 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_428
timestamp 1626908933
transform 1 0 10704 0 1 3071
box -32 -32 32 32
use M1M2_PR  M1M2_PR_892
timestamp 1626908933
transform 1 0 10704 0 1 3515
box -32 -32 32 32
use M1M2_PR  M1M2_PR_427
timestamp 1626908933
transform 1 0 10704 0 1 3515
box -32 -32 32 32
use L1M1_PR  L1M1_PR_559
timestamp 1626908933
transform 1 0 10416 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_57
timestamp 1626908933
transform 1 0 10416 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_522
timestamp 1626908933
transform 1 0 10512 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_57
timestamp 1626908933
transform 1 0 10512 0 1 3663
box -32 -32 32 32
use L1M1_PR  L1M1_PR_971
timestamp 1626908933
transform 1 0 10704 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_743
timestamp 1626908933
transform 1 0 10608 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_469
timestamp 1626908933
transform 1 0 10704 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_241
timestamp 1626908933
transform 1 0 10608 0 1 3663
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_12
timestamp 1626908933
transform 1 0 10272 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_44
timestamp 1626908933
transform 1 0 10272 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_141
timestamp 1626908933
transform 1 0 10944 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_28
timestamp 1626908933
transform 1 0 10944 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_121
timestamp 1626908933
transform 1 0 11136 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_18
timestamp 1626908933
transform 1 0 11136 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_2
timestamp 1626908933
transform 1 0 11904 0 -1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_5
timestamp 1626908933
transform 1 0 11904 0 -1 3996
box -38 -49 518 715
use M1M2_PR  M1M2_PR_102
timestamp 1626908933
transform 1 0 12048 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_103
timestamp 1626908933
transform 1 0 12048 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_567
timestamp 1626908933
transform 1 0 12048 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_568
timestamp 1626908933
transform 1 0 12048 0 1 3219
box -32 -32 32 32
use L1M1_PR  L1M1_PR_98
timestamp 1626908933
transform 1 0 12048 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_426
timestamp 1626908933
transform 1 0 12240 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_600
timestamp 1626908933
transform 1 0 12048 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_928
timestamp 1626908933
transform 1 0 12240 0 1 3663
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_127
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_8
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_127
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_8
timestamp 1626908933
transform 1 0 12500 0 1 3330
box -100 -49 100 49
use L1M1_PR  L1M1_PR_773
timestamp 1626908933
transform 1 0 12432 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_271
timestamp 1626908933
transform 1 0 12432 0 1 3219
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_275
timestamp 1626908933
transform 1 0 12384 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_105
timestamp 1626908933
transform 1 0 12384 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_141
timestamp 1626908933
transform 1 0 12480 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_59
timestamp 1626908933
transform 1 0 12480 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_53
timestamp 1626908933
transform 1 0 12576 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_166
timestamp 1626908933
transform 1 0 12576 0 -1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_220
timestamp 1626908933
transform 1 0 13008 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_221
timestamp 1626908933
transform 1 0 13008 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_685
timestamp 1626908933
transform 1 0 13008 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_686
timestamp 1626908933
transform 1 0 13008 0 1 3219
box -32 -32 32 32
use L1M1_PR  L1M1_PR_775
timestamp 1626908933
transform 1 0 13200 0 1 3219
box -29 -23 29 23
use L1M1_PR  L1M1_PR_273
timestamp 1626908933
transform 1 0 13200 0 1 3219
box -29 -23 29 23
use M1M2_PR  M1M2_PR_688
timestamp 1626908933
transform 1 0 13200 0 1 3219
box -32 -32 32 32
use M1M2_PR  M1M2_PR_223
timestamp 1626908933
transform 1 0 13200 0 1 3219
box -32 -32 32 32
use L1M1_PR  L1M1_PR_774
timestamp 1626908933
transform 1 0 13200 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_772
timestamp 1626908933
transform 1 0 13104 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_272
timestamp 1626908933
transform 1 0 13200 0 1 3663
box -29 -23 29 23
use L1M1_PR  L1M1_PR_270
timestamp 1626908933
transform 1 0 13104 0 1 3663
box -29 -23 29 23
use M1M2_PR  M1M2_PR_842
timestamp 1626908933
transform 1 0 13296 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_687
timestamp 1626908933
transform 1 0 13200 0 1 3663
box -32 -32 32 32
use M1M2_PR  M1M2_PR_377
timestamp 1626908933
transform 1 0 13296 0 1 3441
box -32 -32 32 32
use M1M2_PR  M1M2_PR_222
timestamp 1626908933
transform 1 0 13200 0 1 3663
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_167
timestamp 1626908933
transform 1 0 13440 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_54
timestamp 1626908933
transform 1 0 13440 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_32
timestamp 1626908933
transform -1 0 13440 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_66
timestamp 1626908933
transform -1 0 13440 0 -1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_27
timestamp 1626908933
transform 1 0 13632 0 -1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_56
timestamp 1626908933
transform 1 0 13632 0 -1 3996
box -38 -49 326 715
use M1M2_PR  M1M2_PR_378
timestamp 1626908933
transform 1 0 13680 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_843
timestamp 1626908933
transform 1 0 13680 0 1 3589
box -32 -32 32 32
use L1M1_PR  L1M1_PR_91
timestamp 1626908933
transform 1 0 13680 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_593
timestamp 1626908933
transform 1 0 13680 0 1 3737
box -29 -23 29 23
use M2M3_PR  M2M3_PR_25
timestamp 1626908933
transform 1 0 13680 0 1 3331
box -33 -37 33 37
use M2M3_PR  M2M3_PR_67
timestamp 1626908933
transform 1 0 13680 0 1 3331
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_106
timestamp 1626908933
transform 1 0 13920 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_276
timestamp 1626908933
transform 1 0 13920 0 -1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_376
timestamp 1626908933
transform 1 0 13872 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_841
timestamp 1626908933
transform 1 0 13872 0 1 3737
box -32 -32 32 32
use L1M1_PR  L1M1_PR_424
timestamp 1626908933
transform 1 0 13872 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_926
timestamp 1626908933
transform 1 0 13872 0 1 3737
box -29 -23 29 23
use M1M2_PR  M1M2_PR_844
timestamp 1626908933
transform 1 0 48 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_379
timestamp 1626908933
transform 1 0 48 0 1 4107
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_277
timestamp 1626908933
transform 1 0 192 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_107
timestamp 1626908933
transform 1 0 192 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_140
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_58
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_168
timestamp 1626908933
transform 1 0 0 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_55
timestamp 1626908933
transform 1 0 0 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_236
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_116
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_8
timestamp 1626908933
transform 1 0 912 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_380
timestamp 1626908933
transform 1 0 816 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_473
timestamp 1626908933
transform 1 0 912 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_845
timestamp 1626908933
transform 1 0 816 0 1 3885
box -32 -32 32 32
use L1M1_PR  L1M1_PR_7
timestamp 1626908933
transform 1 0 912 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_509
timestamp 1626908933
transform 1 0 912 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_428
timestamp 1626908933
transform 1 0 1104 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_930
timestamp 1626908933
transform 1 0 1104 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_349
timestamp 1626908933
transform 1 0 1680 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_851
timestamp 1626908933
transform 1 0 1680 0 1 3885
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_116
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_235
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_116
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_235
timestamp 1626908933
transform 1 0 1700 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_218
timestamp 1626908933
transform 1 0 1104 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_683
timestamp 1626908933
transform 1 0 1104 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_459
timestamp 1626908933
transform 1 0 1488 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_924
timestamp 1626908933
transform 1 0 1488 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_42
timestamp 1626908933
transform -1 0 2688 0 1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_5
timestamp 1626908933
transform -1 0 2688 0 1 3996
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_291
timestamp 1626908933
transform 1 0 2256 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_756
timestamp 1626908933
transform 1 0 2256 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_290
timestamp 1626908933
transform 1 0 2256 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_755
timestamp 1626908933
transform 1 0 2256 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_348
timestamp 1626908933
transform 1 0 2256 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_386
timestamp 1626908933
transform 1 0 2736 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_850
timestamp 1626908933
transform 1 0 2256 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_888
timestamp 1626908933
transform 1 0 2736 0 1 4477
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_1
timestamp 1626908933
transform 1 0 2688 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_8
timestamp 1626908933
transform 1 0 2688 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_108
timestamp 1626908933
transform 1 0 3072 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_278
timestamp 1626908933
transform 1 0 3072 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_240
timestamp 1626908933
transform 1 0 2928 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_705
timestamp 1626908933
transform 1 0 2928 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_415
timestamp 1626908933
transform 1 0 3312 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_880
timestamp 1626908933
transform 1 0 3312 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_290
timestamp 1626908933
transform 1 0 3216 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_489
timestamp 1626908933
transform 1 0 3408 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_792
timestamp 1626908933
transform 1 0 3216 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_991
timestamp 1626908933
transform 1 0 3408 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_1
timestamp 1626908933
transform -1 0 3840 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_33
timestamp 1626908933
transform -1 0 3840 0 1 3996
box -38 -49 710 715
use L1M1_PR  L1M1_PR_457
timestamp 1626908933
transform 1 0 3792 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_959
timestamp 1626908933
transform 1 0 3792 0 1 4107
box -29 -23 29 23
use M1M2_PR  M1M2_PR_96
timestamp 1626908933
transform 1 0 3696 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_328
timestamp 1626908933
transform 1 0 3504 0 1 4477
box -32 -32 32 32
use M1M2_PR  M1M2_PR_561
timestamp 1626908933
transform 1 0 3696 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_793
timestamp 1626908933
transform 1 0 3504 0 1 4477
box -32 -32 32 32
use L1M1_PR  L1M1_PR_93
timestamp 1626908933
transform 1 0 3696 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_258
timestamp 1626908933
transform 1 0 3504 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_595
timestamp 1626908933
transform 1 0 3696 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_760
timestamp 1626908933
transform 1 0 3504 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_77
timestamp 1626908933
transform 1 0 3840 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_197
timestamp 1626908933
transform 1 0 3840 0 1 3996
box -38 -49 422 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_225
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_106
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_225
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_106
timestamp 1626908933
transform 1 0 4100 0 1 3996
box -100 -49 100 49
use M1M2_PR  M1M2_PR_758
timestamp 1626908933
transform 1 0 4080 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_293
timestamp 1626908933
transform 1 0 4080 0 1 4551
box -32 -32 32 32
use L1M1_PR  L1M1_PR_852
timestamp 1626908933
transform 1 0 4368 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_350
timestamp 1626908933
transform 1 0 4368 0 1 4551
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_279
timestamp 1626908933
transform 1 0 4224 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_109
timestamp 1626908933
transform 1 0 4224 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_989
timestamp 1626908933
transform 1 0 4560 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_757
timestamp 1626908933
transform 1 0 4656 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_487
timestamp 1626908933
transform 1 0 4560 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_255
timestamp 1626908933
transform 1 0 4656 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_669
timestamp 1626908933
transform 1 0 4656 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_204
timestamp 1626908933
transform 1 0 4656 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_929
timestamp 1626908933
transform 1 0 4944 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_612
timestamp 1626908933
transform 1 0 4944 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_427
timestamp 1626908933
transform 1 0 4944 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_110
timestamp 1626908933
transform 1 0 4944 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_578
timestamp 1626908933
transform 1 0 4944 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_113
timestamp 1626908933
transform 1 0 4944 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_139
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_57
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_31
timestamp 1626908933
transform -1 0 4992 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_63
timestamp 1626908933
transform -1 0 4992 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_68
timestamp 1626908933
transform 1 0 5280 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_188
timestamp 1626908933
transform 1 0 5280 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_27
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_140
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_503
timestamp 1626908933
transform 1 0 5616 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1
timestamp 1626908933
transform 1 0 5616 0 1 3885
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_280
timestamp 1626908933
transform 1 0 5664 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_110
timestamp 1626908933
transform 1 0 5664 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_502
timestamp 1626908933
transform 1 0 5808 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_0
timestamp 1626908933
transform 1 0 5808 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_466
timestamp 1626908933
transform 1 0 5808 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_465
timestamp 1626908933
transform 1 0 5808 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1
timestamp 1626908933
transform 1 0 5808 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_0
timestamp 1626908933
transform 1 0 5808 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__sdlclkp_2  sky130_fd_sc_hs__sdlclkp_2_1
timestamp 1626908933
transform 1 0 5760 0 1 3996
box -38 -49 1670 715
use sky130_fd_sc_hs__sdlclkp_2  sky130_fd_sc_hs__sdlclkp_2_0
timestamp 1626908933
transform 1 0 5760 0 1 3996
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_129
timestamp 1626908933
transform 1 0 6288 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_594
timestamp 1626908933
transform 1 0 6288 0 1 3885
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_96
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_215
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_96
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_215
timestamp 1626908933
transform 1 0 6500 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_133
timestamp 1626908933
transform 1 0 6480 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_635
timestamp 1626908933
transform 1 0 6480 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_285
timestamp 1626908933
transform 1 0 6000 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_787
timestamp 1626908933
transform 1 0 6000 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_200
timestamp 1626908933
transform 1 0 7152 0 1 4181
box -32 -32 32 32
use M1M2_PR  M1M2_PR_436
timestamp 1626908933
transform 1 0 7440 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_665
timestamp 1626908933
transform 1 0 7152 0 1 4181
box -32 -32 32 32
use M1M2_PR  M1M2_PR_901
timestamp 1626908933
transform 1 0 7440 0 1 4107
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1003
timestamp 1626908933
transform 1 0 6864 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_501
timestamp 1626908933
transform 1 0 6864 0 1 4255
box -29 -23 29 23
use M1M2_PR  M1M2_PR_927
timestamp 1626908933
transform 1 0 6864 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_462
timestamp 1626908933
transform 1 0 6864 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_699
timestamp 1626908933
transform 1 0 7056 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_234
timestamp 1626908933
transform 1 0 7056 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_900
timestamp 1626908933
transform 1 0 7440 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_435
timestamp 1626908933
transform 1 0 7440 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_892
timestamp 1626908933
transform 1 0 7248 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_390
timestamp 1626908933
transform 1 0 7248 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_810
timestamp 1626908933
transform 1 0 7440 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_308
timestamp 1626908933
transform 1 0 7440 0 1 4551
box -29 -23 29 23
use M1M2_PR  M1M2_PR_722
timestamp 1626908933
transform 1 0 7440 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_257
timestamp 1626908933
transform 1 0 7440 0 1 4551
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_10
timestamp 1626908933
transform -1 0 8064 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_42
timestamp 1626908933
transform -1 0 8064 0 1 3996
box -38 -49 710 715
use M1M2_PR  M1M2_PR_199
timestamp 1626908933
transform 1 0 7728 0 1 4181
box -32 -32 32 32
use M1M2_PR  M1M2_PR_664
timestamp 1626908933
transform 1 0 7728 0 1 4181
box -32 -32 32 32
use M1M2_PR  M1M2_PR_334
timestamp 1626908933
transform 1 0 7632 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_799
timestamp 1626908933
transform 1 0 7632 0 1 4403
box -32 -32 32 32
use L1M1_PR  L1M1_PR_480
timestamp 1626908933
transform 1 0 7632 0 1 4290
box -29 -23 29 23
use L1M1_PR  L1M1_PR_982
timestamp 1626908933
transform 1 0 7632 0 1 4290
box -29 -23 29 23
use M1M2_PR  M1M2_PR_198
timestamp 1626908933
transform 1 0 7728 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_663
timestamp 1626908933
transform 1 0 7728 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_249
timestamp 1626908933
transform 1 0 7728 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_751
timestamp 1626908933
transform 1 0 7728 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_309
timestamp 1626908933
transform 1 0 7920 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_774
timestamp 1626908933
transform 1 0 7920 0 1 4403
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_86
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_205
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_86
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_205
timestamp 1626908933
transform 1 0 8900 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_448
timestamp 1626908933
transform 1 0 8016 0 1 4107
box -29 -23 29 23
use L1M1_PR  L1M1_PR_950
timestamp 1626908933
transform 1 0 8016 0 1 4107
box -29 -23 29 23
use M1M2_PR  M1M2_PR_406
timestamp 1626908933
transform 1 0 8592 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_871
timestamp 1626908933
transform 1 0 8592 0 1 4107
box -32 -32 32 32
use M1M2_PR  M1M2_PR_65
timestamp 1626908933
transform 1 0 8016 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_530
timestamp 1626908933
transform 1 0 8016 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_64
timestamp 1626908933
transform 1 0 8016 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_566
timestamp 1626908933
transform 1 0 8016 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_333
timestamp 1626908933
transform 1 0 8400 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_798
timestamp 1626908933
transform 1 0 8400 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_389
timestamp 1626908933
transform 1 0 8400 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_891
timestamp 1626908933
transform 1 0 8400 0 1 4329
box -29 -23 29 23
use M2M3_PR  M2M3_PR_3
timestamp 1626908933
transform 1 0 8016 0 1 4551
box -33 -37 33 37
use M2M3_PR  M2M3_PR_45
timestamp 1626908933
transform 1 0 8016 0 1 4551
box -33 -37 33 37
use M1M2_PR  M1M2_PR_149
timestamp 1626908933
transform 1 0 8304 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_614
timestamp 1626908933
transform 1 0 8304 0 1 4551
box -32 -32 32 32
use M2M3_PR  M2M3_PR_2
timestamp 1626908933
transform 1 0 8400 0 1 4551
box -33 -37 33 37
use M2M3_PR  M2M3_PR_44
timestamp 1626908933
transform 1 0 8400 0 1 4551
box -33 -37 33 37
use M1M2_PR  M1M2_PR_258
timestamp 1626908933
transform 1 0 9072 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_308
timestamp 1626908933
transform 1 0 9072 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_723
timestamp 1626908933
transform 1 0 9072 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_773
timestamp 1626908933
transform 1 0 9072 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_405
timestamp 1626908933
transform 1 0 9360 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_870
timestamp 1626908933
transform 1 0 9360 0 1 3811
box -32 -32 32 32
use L1M1_PR  L1M1_PR_310
timestamp 1626908933
transform 1 0 9552 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_812
timestamp 1626908933
transform 1 0 9552 0 1 3885
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_56
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_138
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_81
timestamp 1626908933
transform 1 0 9936 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_546
timestamp 1626908933
transform 1 0 9936 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_16  sky130_fd_sc_hs__clkbuf_16_0
timestamp 1626908933
transform 1 0 8064 0 1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  sky130_fd_sc_hs__clkbuf_16_1
timestamp 1626908933
transform 1 0 8064 0 1 3996
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_949
timestamp 1626908933
transform 1 0 10128 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_447
timestamp 1626908933
transform 1 0 10128 0 1 3885
box -29 -23 29 23
use M1M2_PR  M1M2_PR_894
timestamp 1626908933
transform 1 0 10128 0 1 4181
box -32 -32 32 32
use M1M2_PR  M1M2_PR_429
timestamp 1626908933
transform 1 0 10128 0 1 4181
box -32 -32 32 32
use L1M1_PR  L1M1_PR_948
timestamp 1626908933
transform 1 0 10320 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_564
timestamp 1626908933
transform 1 0 10224 0 1 3811
box -29 -23 29 23
use L1M1_PR  L1M1_PR_446
timestamp 1626908933
transform 1 0 10320 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_62
timestamp 1626908933
transform 1 0 10224 0 1 3811
box -29 -23 29 23
use M1M2_PR  M1M2_PR_768
timestamp 1626908933
transform 1 0 10320 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_303
timestamp 1626908933
transform 1 0 10320 0 1 4403
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_234
timestamp 1626908933
transform 1 0 10272 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_64
timestamp 1626908933
transform 1 0 10272 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_139
timestamp 1626908933
transform 1 0 10080 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_26
timestamp 1626908933
transform 1 0 10080 0 1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_61
timestamp 1626908933
transform 1 0 10704 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_404
timestamp 1626908933
transform 1 0 10416 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_526
timestamp 1626908933
transform 1 0 10704 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_869
timestamp 1626908933
transform 1 0 10416 0 1 3885
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_25
timestamp 1626908933
transform 1 0 10368 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_128
timestamp 1626908933
transform 1 0 10368 0 1 3996
box -38 -49 806 715
use M1M2_PR  M1M2_PR_261
timestamp 1626908933
transform 1 0 11088 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_726
timestamp 1626908933
transform 1 0 11088 0 1 3885
box -32 -32 32 32
use L1M1_PR  L1M1_PR_313
timestamp 1626908933
transform 1 0 10896 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_815
timestamp 1626908933
transform 1 0 10896 0 1 3885
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_76
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_195
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_76
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_195
timestamp 1626908933
transform 1 0 11300 0 1 3996
box -100 -49 100 49
use L1M1_PR  L1M1_PR_922
timestamp 1626908933
transform 1 0 11472 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_729
timestamp 1626908933
transform 1 0 11280 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_581
timestamp 1626908933
transform 1 0 11280 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_420
timestamp 1626908933
transform 1 0 11472 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_227
timestamp 1626908933
transform 1 0 11280 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_79
timestamp 1626908933
transform 1 0 11280 0 1 4329
box -29 -23 29 23
use M1M2_PR  M1M2_PR_647
timestamp 1626908933
transform 1 0 11280 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_182
timestamp 1626908933
transform 1 0 11280 0 1 4551
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_138
timestamp 1626908933
transform 1 0 11616 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_25
timestamp 1626908933
transform 1 0 11616 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_4
timestamp 1626908933
transform 1 0 11136 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_1
timestamp 1626908933
transform 1 0 11136 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_233
timestamp 1626908933
transform 1 0 11808 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_63
timestamp 1626908933
transform 1 0 11808 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_137
timestamp 1626908933
transform 1 0 11904 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_17
timestamp 1626908933
transform 1 0 11904 0 1 3996
box -38 -49 422 715
use M1M2_PR  M1M2_PR_181
timestamp 1626908933
transform 1 0 12048 0 1 3811
box -32 -32 32 32
use M1M2_PR  M1M2_PR_646
timestamp 1626908933
transform 1 0 12048 0 1 3811
box -32 -32 32 32
use L1M1_PR  L1M1_PR_225
timestamp 1626908933
transform 1 0 12240 0 1 3811
box -29 -23 29 23
use L1M1_PR  L1M1_PR_727
timestamp 1626908933
transform 1 0 12240 0 1 3811
box -29 -23 29 23
use M1M2_PR  M1M2_PR_233
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_698
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -32 -32 32 32
use L1M1_PR  L1M1_PR_282
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_287
timestamp 1626908933
transform 1 0 12720 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_465
timestamp 1626908933
transform 1 0 12528 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_784
timestamp 1626908933
transform 1 0 12336 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_789
timestamp 1626908933
transform 1 0 12720 0 1 4255
box -29 -23 29 23
use L1M1_PR  L1M1_PR_967
timestamp 1626908933
transform 1 0 12528 0 1 4255
box -29 -23 29 23
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_5
timestamp 1626908933
transform -1 0 12768 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__nor2b_1  sky130_fd_sc_hs__nor2b_1_11
timestamp 1626908933
transform -1 0 12768 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_56
timestamp 1626908933
transform 1 0 12768 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_169
timestamp 1626908933
transform 1 0 12768 0 1 3996
box -38 -49 230 715
use L1M1_PR  L1M1_PR_286
timestamp 1626908933
transform 1 0 12816 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_788
timestamp 1626908933
transform 1 0 12816 0 1 3885
box -29 -23 29 23
use M1M2_PR  M1M2_PR_702
timestamp 1626908933
transform 1 0 13104 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_237
timestamp 1626908933
transform 1 0 13104 0 1 3885
box -32 -32 32 32
use M2M3_PR  M2M3_PR_66
timestamp 1626908933
transform 1 0 13296 0 1 3941
box -33 -37 33 37
use M2M3_PR  M2M3_PR_24
timestamp 1626908933
transform 1 0 13296 0 1 3941
box -33 -37 33 37
use M1M2_PR  M1M2_PR_835
timestamp 1626908933
transform 1 0 13200 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_701
timestamp 1626908933
transform 1 0 13104 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_370
timestamp 1626908933
transform 1 0 13200 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_236
timestamp 1626908933
transform 1 0 13104 0 1 4255
box -32 -32 32 32
use L1M1_PR  L1M1_PR_894
timestamp 1626908933
transform 1 0 13296 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_392
timestamp 1626908933
transform 1 0 13296 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_663
timestamp 1626908933
transform 1 0 13200 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_161
timestamp 1626908933
transform 1 0 13200 0 1 4477
box -29 -23 29 23
use L1M1_PR  L1M1_PR_666
timestamp 1626908933
transform 1 0 13296 0 1 4403
box -29 -23 29 23
use L1M1_PR  L1M1_PR_164
timestamp 1626908933
transform 1 0 13296 0 1 4403
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_13
timestamp 1626908933
transform -1 0 13632 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_47
timestamp 1626908933
transform -1 0 13632 0 1 3996
box -38 -49 710 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_55
timestamp 1626908933
transform 1 0 13632 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_137
timestamp 1626908933
transform 1 0 13632 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_57
timestamp 1626908933
transform 1 0 13728 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_170
timestamp 1626908933
transform 1 0 13728 0 1 3996
box -38 -49 230 715
use M1M2_PR  M1M2_PR_151
timestamp 1626908933
transform 1 0 13680 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_336
timestamp 1626908933
transform 1 0 13488 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_616
timestamp 1626908933
transform 1 0 13680 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_801
timestamp 1626908933
transform 1 0 13488 0 1 4329
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_111
timestamp 1626908933
transform 1 0 13920 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_281
timestamp 1626908933
transform 1 0 13920 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_189
timestamp 1626908933
transform 1 0 13968 0 1 3885
box -32 -32 32 32
use M1M2_PR  M1M2_PR_654
timestamp 1626908933
transform 1 0 13968 0 1 3885
box -32 -32 32 32
use L1M1_PR  L1M1_PR_235
timestamp 1626908933
transform 1 0 13872 0 1 3885
box -29 -23 29 23
use L1M1_PR  L1M1_PR_737
timestamp 1626908933
transform 1 0 13872 0 1 3885
box -29 -23 29 23
use M2M3_PR  M2M3_PR_23
timestamp 1626908933
transform 1 0 13776 0 1 4551
box -33 -37 33 37
use M2M3_PR  M2M3_PR_65
timestamp 1626908933
transform 1 0 13776 0 1 4551
box -33 -37 33 37
use M2M3_PR  M2M3_PR_72
timestamp 1626908933
transform 1 0 48 0 1 4795
box -33 -37 33 37
use M2M3_PR  M2M3_PR_30
timestamp 1626908933
transform 1 0 48 0 1 4795
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_284
timestamp 1626908933
transform 1 0 192 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_114
timestamp 1626908933
transform 1 0 192 0 1 5328
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_181
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_62
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_181
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_62
timestamp 1626908933
transform 1 0 500 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_133
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_51
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_175
timestamp 1626908933
transform 1 0 0 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_62
timestamp 1626908933
transform 1 0 0 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_235
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_115
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_7
timestamp 1626908933
transform 1 0 912 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_381
timestamp 1626908933
transform 1 0 720 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_472
timestamp 1626908933
transform 1 0 912 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_846
timestamp 1626908933
transform 1 0 720 0 1 5217
box -32 -32 32 32
use L1M1_PR  L1M1_PR_6
timestamp 1626908933
transform 1 0 912 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_429
timestamp 1626908933
transform 1 0 816 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_508
timestamp 1626908933
transform 1 0 912 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_931
timestamp 1626908933
transform 1 0 816 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_89
timestamp 1626908933
transform 1 0 768 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_99
timestamp 1626908933
transform 1 0 0 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_192
timestamp 1626908933
transform 1 0 768 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_202
timestamp 1626908933
transform 1 0 0 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_29
timestamp 1626908933
transform 1 0 768 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_61
timestamp 1626908933
transform 1 0 768 0 -1 5328
box -38 -49 710 715
use M1M2_PR  M1M2_PR_469
timestamp 1626908933
transform 1 0 1296 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_4
timestamp 1626908933
transform 1 0 1296 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_217
timestamp 1626908933
transform 1 0 1104 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_682
timestamp 1626908933
transform 1 0 1104 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_269
timestamp 1626908933
transform 1 0 1104 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_771
timestamp 1626908933
transform 1 0 1104 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_500
timestamp 1626908933
transform 1 0 1200 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1002
timestamp 1626908933
transform 1 0 1200 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_458
timestamp 1626908933
transform 1 0 1488 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_923
timestamp 1626908933
transform 1 0 1488 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_289
timestamp 1626908933
transform 1 0 1392 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_754
timestamp 1626908933
transform 1 0 1392 0 1 5217
box -32 -32 32 32
use L1M1_PR  L1M1_PR_347
timestamp 1626908933
transform 1 0 1392 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_849
timestamp 1626908933
transform 1 0 1392 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_137
timestamp 1626908933
transform 1 0 1440 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_24
timestamp 1626908933
transform 1 0 1440 0 -1 5328
box -38 -49 230 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_234
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_115
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_234
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_115
timestamp 1626908933
transform 1 0 1700 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_232
timestamp 1626908933
transform 1 0 1632 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_62
timestamp 1626908933
transform 1 0 1632 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_920
timestamp 1626908933
transform 1 0 1968 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_455
timestamp 1626908933
transform 1 0 1968 0 1 4995
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_221
timestamp 1626908933
transform 1 0 1536 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_101
timestamp 1626908933
transform 1 0 1536 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_75
timestamp 1626908933
transform 1 0 1728 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_178
timestamp 1626908933
transform 1 0 1728 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_67
timestamp 1626908933
transform -1 0 3840 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_30
timestamp 1626908933
transform -1 0 3840 0 1 5328
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_170
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_51
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_170
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_51
timestamp 1626908933
transform 1 0 2900 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_505
timestamp 1626908933
transform 1 0 2736 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3
timestamp 1626908933
transform 1 0 2736 0 1 4773
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_136
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_54
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_792
timestamp 1626908933
transform 1 0 3504 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_468
timestamp 1626908933
transform 1 0 3888 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_327
timestamp 1626908933
transform 1 0 3504 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3
timestamp 1626908933
transform 1 0 3888 0 1 4773
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_196
timestamp 1626908933
transform 1 0 3840 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_76
timestamp 1626908933
transform 1 0 3840 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_68
timestamp 1626908933
transform -1 0 4512 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_31
timestamp 1626908933
transform -1 0 4512 0 -1 5328
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_224
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_105
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_224
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_105
timestamp 1626908933
transform 1 0 4100 0 1 5328
box -100 -49 100 49
use L1M1_PR  L1M1_PR_853
timestamp 1626908933
transform 1 0 4080 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_351
timestamp 1626908933
transform 1 0 4080 0 1 5069
box -29 -23 29 23
use M1M2_PR  M1M2_PR_757
timestamp 1626908933
transform 1 0 4080 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_292
timestamp 1626908933
transform 1 0 4080 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_285
timestamp 1626908933
transform 1 0 4416 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_115
timestamp 1626908933
transform 1 0 4416 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_176
timestamp 1626908933
transform 1 0 4224 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_63
timestamp 1626908933
transform 1 0 4224 0 1 5328
box -38 -49 230 715
use L1M1_PR  L1M1_PR_878
timestamp 1626908933
transform 1 0 4464 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_376
timestamp 1626908933
transform 1 0 4464 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_282
timestamp 1626908933
transform 1 0 4896 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_112
timestamp 1626908933
transform 1 0 4896 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_177
timestamp 1626908933
transform 1 0 4800 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_64
timestamp 1626908933
transform 1 0 4800 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_193
timestamp 1626908933
transform 1 0 4512 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_73
timestamp 1626908933
transform 1 0 4512 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_40
timestamp 1626908933
transform 1 0 4512 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_11
timestamp 1626908933
transform 1 0 4512 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_50
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_132
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_309
timestamp 1626908933
transform 1 0 5424 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_375
timestamp 1626908933
transform 1 0 5040 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_811
timestamp 1626908933
transform 1 0 5424 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_877
timestamp 1626908933
transform 1 0 5040 0 1 4995
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_40
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_159
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_40
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_159
timestamp 1626908933
transform 1 0 5300 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_2
timestamp 1626908933
transform 1 0 5760 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_9
timestamp 1626908933
transform 1 0 5760 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_15
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_49
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_52
timestamp 1626908933
transform 1 0 4992 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_15
timestamp 1626908933
transform 1 0 4992 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_14
timestamp 1626908933
transform 1 0 6144 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_43
timestamp 1626908933
transform 1 0 6144 0 1 5328
box -38 -49 326 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_95
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_214
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_95
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_214
timestamp 1626908933
transform 1 0 6500 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_23
timestamp 1626908933
transform 1 0 6912 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_136
timestamp 1626908933
transform 1 0 6912 0 -1 5328
box -38 -49 230 715
use L1M1_PR  L1M1_PR_68
timestamp 1626908933
transform 1 0 6768 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_570
timestamp 1626908933
transform 1 0 6768 0 1 4773
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_19
timestamp 1626908933
transform 1 0 6432 0 1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_53
timestamp 1626908933
transform 1 0 6432 0 1 5328
box -38 -49 710 715
use M1M2_PR  M1M2_PR_721
timestamp 1626908933
transform 1 0 7440 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_532
timestamp 1626908933
transform 1 0 7248 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_256
timestamp 1626908933
transform 1 0 7440 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_67
timestamp 1626908933
transform 1 0 7248 0 1 4773
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_135
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_53
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_177
timestamp 1626908933
transform 1 0 7104 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_57
timestamp 1626908933
transform 1 0 7104 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_44
timestamp 1626908933
transform 1 0 7104 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_15
timestamp 1626908933
transform 1 0 7104 0 1 5328
box -38 -49 326 715
use L1M1_PR  L1M1_PR_65
timestamp 1626908933
transform 1 0 7920 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_567
timestamp 1626908933
transform 1 0 7920 0 1 5143
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_29
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_148
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_29
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_148
timestamp 1626908933
transform 1 0 7700 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_12
timestamp 1626908933
transform 1 0 7392 0 1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_46
timestamp 1626908933
transform 1 0 7392 0 1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_53
timestamp 1626908933
transform -1 0 9504 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_16
timestamp 1626908933
transform -1 0 9504 0 -1 5328
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_204
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_85
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_204
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_85
timestamp 1626908933
transform 1 0 8900 0 1 5328
box -100 -49 100 49
use M1M2_PR  M1M2_PR_724
timestamp 1626908933
transform 1 0 8880 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_529
timestamp 1626908933
transform 1 0 8112 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_259
timestamp 1626908933
transform 1 0 8880 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_64
timestamp 1626908933
transform 1 0 8112 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_307
timestamp 1626908933
transform 1 0 9072 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_772
timestamp 1626908933
transform 1 0 9072 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_311
timestamp 1626908933
transform 1 0 9088 0 1 4884
box -29 -23 29 23
use L1M1_PR  L1M1_PR_364
timestamp 1626908933
transform 1 0 9456 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_813
timestamp 1626908933
transform 1 0 9088 0 1 4884
box -29 -23 29 23
use L1M1_PR  L1M1_PR_866
timestamp 1626908933
transform 1 0 9456 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_728
timestamp 1626908933
transform 1 0 9648 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_263
timestamp 1626908933
transform 1 0 9648 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_194
timestamp 1626908933
transform 1 0 9744 0 1 4847
box -32 -32 32 32
use M1M2_PR  M1M2_PR_659
timestamp 1626908933
transform 1 0 9744 0 1 4847
box -32 -32 32 32
use M1M2_PR  M1M2_PR_63
timestamp 1626908933
transform 1 0 9936 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_431
timestamp 1626908933
transform 1 0 9936 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_528
timestamp 1626908933
transform 1 0 9936 0 1 5143
box -32 -32 32 32
use M1M2_PR  M1M2_PR_896
timestamp 1626908933
transform 1 0 9936 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_314
timestamp 1626908933
transform 1 0 9744 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_471
timestamp 1626908933
transform 1 0 9936 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_816
timestamp 1626908933
transform 1 0 9744 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_973
timestamp 1626908933
transform 1 0 9936 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_49
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_131
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_171
timestamp 1626908933
transform 1 0 9504 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_58
timestamp 1626908933
transform 1 0 9504 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_13
timestamp 1626908933
transform -1 0 10368 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_45
timestamp 1626908933
transform -1 0 10368 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_39
timestamp 1626908933
transform -1 0 9984 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_2
timestamp 1626908933
transform -1 0 9984 0 1 5328
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_137
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_18
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_137
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_18
timestamp 1626908933
transform 1 0 10100 0 1 4662
box -100 -49 100 49
use L1M1_PR  L1M1_PR_242
timestamp 1626908933
transform 1 0 10032 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_744
timestamp 1626908933
transform 1 0 10032 0 1 4995
box -29 -23 29 23
use M1M2_PR  M1M2_PR_302
timestamp 1626908933
transform 1 0 10320 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_767
timestamp 1626908933
transform 1 0 10320 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_445
timestamp 1626908933
transform 1 0 10320 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_947
timestamp 1626908933
transform 1 0 10320 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_55
timestamp 1626908933
transform 1 0 10416 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_557
timestamp 1626908933
transform 1 0 10416 0 1 5217
box -29 -23 29 23
use M2M3_PR  M2M3_PR_1
timestamp 1626908933
transform 1 0 10320 0 1 5283
box -33 -37 33 37
use M2M3_PR  M2M3_PR_43
timestamp 1626908933
transform 1 0 10320 0 1 5283
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_172
timestamp 1626908933
transform 1 0 10368 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_59
timestamp 1626908933
transform 1 0 10368 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_155
timestamp 1626908933
transform 1 0 10080 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_35
timestamp 1626908933
transform 1 0 10080 0 1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_55
timestamp 1626908933
transform 1 0 10704 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_60
timestamp 1626908933
transform 1 0 10704 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_403
timestamp 1626908933
transform 1 0 10800 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_520
timestamp 1626908933
transform 1 0 10704 0 1 5217
box -32 -32 32 32
use M1M2_PR  M1M2_PR_525
timestamp 1626908933
transform 1 0 10704 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_868
timestamp 1626908933
transform 1 0 10800 0 1 5069
box -32 -32 32 32
use L1M1_PR  L1M1_PR_359
timestamp 1626908933
transform 1 0 10608 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_861
timestamp 1626908933
transform 1 0 10608 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_24
timestamp 1626908933
transform 1 0 10464 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_127
timestamp 1626908933
transform 1 0 10464 0 1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_260
timestamp 1626908933
transform 1 0 11088 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_725
timestamp 1626908933
transform 1 0 11088 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_312
timestamp 1626908933
transform 1 0 10992 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_814
timestamp 1626908933
transform 1 0 10992 0 1 4995
box -29 -23 29 23
use M2M3_PR  M2M3_PR_0
timestamp 1626908933
transform 1 0 11088 0 1 5283
box -33 -37 33 37
use M2M3_PR  M2M3_PR_42
timestamp 1626908933
transform 1 0 11088 0 1 5283
box -33 -37 33 37
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_75
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_194
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_75
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_194
timestamp 1626908933
transform 1 0 11300 0 1 5328
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_178
timestamp 1626908933
transform 1 0 11232 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_65
timestamp 1626908933
transform 1 0 11232 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_73
timestamp 1626908933
transform 1 0 11424 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_38
timestamp 1626908933
transform 1 0 10560 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_36
timestamp 1626908933
transform 1 0 11424 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_1
timestamp 1626908933
transform 1 0 10560 0 -1 5328
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_61
timestamp 1626908933
transform 1 0 12144 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_563
timestamp 1626908933
transform 1 0 12144 0 1 4773
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_52
timestamp 1626908933
transform 1 0 12480 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_134
timestamp 1626908933
transform 1 0 12480 0 -1 5328
box -38 -49 134 715
use L1M1_PR  L1M1_PR_60
timestamp 1626908933
transform 1 0 12336 0 1 5143
box -29 -23 29 23
use L1M1_PR  L1M1_PR_562
timestamp 1626908933
transform 1 0 12336 0 1 5143
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_7
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_126
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_7
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_126
timestamp 1626908933
transform 1 0 12500 0 1 4662
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_60
timestamp 1626908933
transform 1 0 12576 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_173
timestamp 1626908933
transform 1 0 12576 0 -1 5328
box -38 -49 230 715
use L1M1_PR  L1M1_PR_916
timestamp 1626908933
transform 1 0 13008 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_670
timestamp 1626908933
transform 1 0 12912 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_561
timestamp 1626908933
transform 1 0 12816 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_414
timestamp 1626908933
transform 1 0 13008 0 1 5069
box -29 -23 29 23
use L1M1_PR  L1M1_PR_168
timestamp 1626908933
transform 1 0 12912 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_59
timestamp 1626908933
transform 1 0 12816 0 1 5069
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_174
timestamp 1626908933
transform 1 0 13056 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_61
timestamp 1626908933
transform 1 0 13056 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_37
timestamp 1626908933
transform 1 0 12768 0 -1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_8
timestamp 1626908933
transform 1 0 12768 0 -1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_66
timestamp 1626908933
transform 1 0 13344 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_179
timestamp 1626908933
transform 1 0 13344 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_113
timestamp 1626908933
transform 1 0 13248 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_283
timestamp 1626908933
transform 1 0 13248 0 -1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_360
timestamp 1626908933
transform 1 0 13200 0 1 5069
box -32 -32 32 32
use M1M2_PR  M1M2_PR_825
timestamp 1626908933
transform 1 0 13200 0 1 5069
box -32 -32 32 32
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_14
timestamp 1626908933
transform 1 0 13344 0 -1 5328
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_48
timestamp 1626908933
transform 1 0 13344 0 -1 5328
box -38 -49 710 715
use M1M2_PR  M1M2_PR_615
timestamp 1626908933
transform 1 0 13680 0 1 4773
box -32 -32 32 32
use M1M2_PR  M1M2_PR_150
timestamp 1626908933
transform 1 0 13680 0 1 4773
box -32 -32 32 32
use M2M3_PR  M2M3_PR_64
timestamp 1626908933
transform 1 0 13584 0 1 5283
box -33 -37 33 37
use M2M3_PR  M2M3_PR_22
timestamp 1626908933
transform 1 0 13584 0 1 5283
box -33 -37 33 37
use L1M1_PR  L1M1_PR_669
timestamp 1626908933
transform 1 0 13584 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_668
timestamp 1626908933
transform 1 0 13680 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_167
timestamp 1626908933
transform 1 0 13584 0 1 4995
box -29 -23 29 23
use L1M1_PR  L1M1_PR_166
timestamp 1626908933
transform 1 0 13680 0 1 4995
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_286
timestamp 1626908933
transform 1 0 13536 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_116
timestamp 1626908933
transform 1 0 13536 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_180
timestamp 1626908933
transform 1 0 13728 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_67
timestamp 1626908933
transform 1 0 13728 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_130
timestamp 1626908933
transform 1 0 13632 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_48
timestamp 1626908933
transform 1 0 13632 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_117
timestamp 1626908933
transform 1 0 13920 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_287
timestamp 1626908933
transform 1 0 13920 0 1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_153
timestamp 1626908933
transform 1 0 13776 0 1 4995
box -32 -32 32 32
use M1M2_PR  M1M2_PR_618
timestamp 1626908933
transform 1 0 13776 0 1 4995
box -32 -32 32 32
use L1M1_PR  L1M1_PR_163
timestamp 1626908933
transform 1 0 13776 0 1 4773
box -29 -23 29 23
use L1M1_PR  L1M1_PR_665
timestamp 1626908933
transform 1 0 13776 0 1 4773
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_180
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_61
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_180
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_61
timestamp 1626908933
transform 1 0 500 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_231
timestamp 1626908933
transform 1 0 0 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_61
timestamp 1626908933
transform 1 0 0 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_201
timestamp 1626908933
transform 1 0 96 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_98
timestamp 1626908933
transform 1 0 96 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_10
timestamp 1626908933
transform 1 0 960 0 -1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_39
timestamp 1626908933
transform 1 0 960 0 -1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_68
timestamp 1626908933
transform 1 0 1248 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_181
timestamp 1626908933
transform 1 0 1248 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_60
timestamp 1626908933
transform 1 0 864 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_230
timestamp 1626908933
transform 1 0 864 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_118
timestamp 1626908933
transform 1 0 1440 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_288
timestamp 1626908933
transform 1 0 1440 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_288
timestamp 1626908933
transform 1 0 1392 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_753
timestamp 1626908933
transform 1 0 1392 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_28
timestamp 1626908933
transform 1 0 1536 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_60
timestamp 1626908933
transform 1 0 1536 0 -1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_477
timestamp 1626908933
transform 1 0 1776 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_12
timestamp 1626908933
transform 1 0 1776 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_69
timestamp 1626908933
transform 1 0 2208 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_182
timestamp 1626908933
transform 1 0 2208 0 -1 6660
box -38 -49 230 715
use L1M1_PR  L1M1_PR_9
timestamp 1626908933
transform 1 0 2064 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_511
timestamp 1626908933
transform 1 0 2064 0 1 5883
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_47
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_129
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_119
timestamp 1626908933
transform 1 0 2400 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_289
timestamp 1626908933
transform 1 0 2400 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_10
timestamp 1626908933
transform 1 0 2352 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_475
timestamp 1626908933
transform 1 0 2352 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_70
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_183
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_155
timestamp 1626908933
transform 1 0 2736 0 1 5809
box -32 -32 32 32
use M1M2_PR  M1M2_PR_620
timestamp 1626908933
transform 1 0 2736 0 1 5809
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_50
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_169
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_50
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_169
timestamp 1626908933
transform 1 0 2900 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_881
timestamp 1626908933
transform 1 0 3792 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_848
timestamp 1626908933
transform 1 0 3408 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_379
timestamp 1626908933
transform 1 0 3792 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_346
timestamp 1626908933
transform 1 0 3408 0 1 5587
box -29 -23 29 23
use M1M2_PR  M1M2_PR_791
timestamp 1626908933
transform 1 0 3504 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_556
timestamp 1626908933
transform 1 0 3696 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_326
timestamp 1626908933
transform 1 0 3504 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_91
timestamp 1626908933
transform 1 0 3696 0 1 5587
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_41
timestamp 1626908933
transform 1 0 2784 0 -1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_4
timestamp 1626908933
transform 1 0 2784 0 -1 6660
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_672
timestamp 1626908933
transform 1 0 4656 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_587
timestamp 1626908933
transform 1 0 4560 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_170
timestamp 1626908933
transform 1 0 4656 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_85
timestamp 1626908933
transform 1 0 4560 0 1 5587
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_157
timestamp 1626908933
transform 1 0 4704 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_54
timestamp 1626908933
transform 1 0 4704 0 -1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_169
timestamp 1626908933
transform 1 0 5424 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_422
timestamp 1626908933
transform 1 0 4848 0 1 5513
box -29 -23 29 23
use L1M1_PR  L1M1_PR_671
timestamp 1626908933
transform 1 0 5424 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_924
timestamp 1626908933
transform 1 0 4848 0 1 5513
box -29 -23 29 23
use L1M1_PR  L1M1_PR_160
timestamp 1626908933
transform 1 0 5520 0 1 5809
box -29 -23 29 23
use L1M1_PR  L1M1_PR_171
timestamp 1626908933
transform 1 0 5424 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_662
timestamp 1626908933
transform 1 0 5520 0 1 5809
box -29 -23 29 23
use L1M1_PR  L1M1_PR_673
timestamp 1626908933
transform 1 0 5424 0 1 5735
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_39
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_158
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_39
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_158
timestamp 1626908933
transform 1 0 5300 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_5
timestamp 1626908933
transform 1 0 5472 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_39
timestamp 1626908933
transform 1 0 5472 0 -1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_70
timestamp 1626908933
transform 1 0 6000 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_92
timestamp 1626908933
transform 1 0 6672 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_535
timestamp 1626908933
transform 1 0 6000 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_557
timestamp 1626908933
transform 1 0 6672 0 1 5513
box -32 -32 32 32
use L1M1_PR  L1M1_PR_70
timestamp 1626908933
transform 1 0 6096 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_417
timestamp 1626908933
transform 1 0 6384 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_572
timestamp 1626908933
transform 1 0 6096 0 1 5439
box -29 -23 29 23
use L1M1_PR  L1M1_PR_919
timestamp 1626908933
transform 1 0 6384 0 1 5587
box -29 -23 29 23
use M1M2_PR  M1M2_PR_160
timestamp 1626908933
transform 1 0 6480 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_625
timestamp 1626908933
transform 1 0 6480 0 1 5883
box -32 -32 32 32
use L1M1_PR  L1M1_PR_188
timestamp 1626908933
transform 1 0 6288 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_690
timestamp 1626908933
transform 1 0 6288 0 1 5735
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_18
timestamp 1626908933
transform 1 0 6144 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_52
timestamp 1626908933
transform 1 0 6144 0 -1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_367
timestamp 1626908933
transform 1 0 6864 0 1 5587
box -32 -32 32 32
use M1M2_PR  M1M2_PR_832
timestamp 1626908933
transform 1 0 6864 0 1 5587
box -32 -32 32 32
use L1M1_PR  L1M1_PR_183
timestamp 1626908933
transform 1 0 6864 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_186
timestamp 1626908933
transform 1 0 6768 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_187
timestamp 1626908933
transform 1 0 6768 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_685
timestamp 1626908933
transform 1 0 6864 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_688
timestamp 1626908933
transform 1 0 6768 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_689
timestamp 1626908933
transform 1 0 6768 0 1 5735
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_46
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_128
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_88
timestamp 1626908933
transform 1 0 7152 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_185
timestamp 1626908933
transform 1 0 7248 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_423
timestamp 1626908933
transform 1 0 7344 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_590
timestamp 1626908933
transform 1 0 7152 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_687
timestamp 1626908933
transform 1 0 7248 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_925
timestamp 1626908933
transform 1 0 7344 0 1 5587
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_17
timestamp 1626908933
transform 1 0 6816 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_51
timestamp 1626908933
transform 1 0 6816 0 -1 6660
box -38 -49 710 715
use L1M1_PR  L1M1_PR_661
timestamp 1626908933
transform 1 0 7728 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_159
timestamp 1626908933
transform 1 0 7728 0 1 5661
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_147
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_28
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_147
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_28
timestamp 1626908933
transform 1 0 7700 0 1 5994
box -100 -49 100 49
use L1M1_PR  L1M1_PR_664
timestamp 1626908933
transform 1 0 7728 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_654
timestamp 1626908933
transform 1 0 7824 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_162
timestamp 1626908933
transform 1 0 7728 0 1 5735
box -29 -23 29 23
use L1M1_PR  L1M1_PR_152
timestamp 1626908933
transform 1 0 7824 0 1 5883
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_229
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_59
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_53
timestamp 1626908933
transform 1 0 7680 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_173
timestamp 1626908933
transform 1 0 7680 0 -1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_59
timestamp 1626908933
transform 1 0 8400 0 1 5809
box -32 -32 32 32
use M1M2_PR  M1M2_PR_148
timestamp 1626908933
transform 1 0 8304 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_524
timestamp 1626908933
transform 1 0 8400 0 1 5809
box -32 -32 32 32
use M1M2_PR  M1M2_PR_613
timestamp 1626908933
transform 1 0 8304 0 1 5735
box -32 -32 32 32
use L1M1_PR  L1M1_PR_58
timestamp 1626908933
transform 1 0 8400 0 1 5809
box -29 -23 29 23
use L1M1_PR  L1M1_PR_560
timestamp 1626908933
transform 1 0 8400 0 1 5809
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_58
timestamp 1626908933
transform 1 0 8832 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_228
timestamp 1626908933
transform 1 0 8832 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_373
timestamp 1626908933
transform 1 0 8496 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_374
timestamp 1626908933
transform 1 0 8496 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_838
timestamp 1626908933
transform 1 0 8496 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_839
timestamp 1626908933
transform 1 0 8496 0 1 5439
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_35
timestamp 1626908933
transform 1 0 8064 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_138
timestamp 1626908933
transform 1 0 8064 0 -1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_262
timestamp 1626908933
transform 1 0 9648 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_306
timestamp 1626908933
transform 1 0 9072 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_727
timestamp 1626908933
transform 1 0 9648 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_771
timestamp 1626908933
transform 1 0 9072 0 1 5661
box -32 -32 32 32
use L1M1_PR  L1M1_PR_315
timestamp 1626908933
transform 1 0 9552 0 1 5587
box -29 -23 29 23
use L1M1_PR  L1M1_PR_817
timestamp 1626908933
transform 1 0 9552 0 1 5587
box -29 -23 29 23
use M1M2_PR  M1M2_PR_141
timestamp 1626908933
transform 1 0 9072 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_606
timestamp 1626908933
transform 1 0 9072 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_29
timestamp 1626908933
transform 1 0 9312 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_132
timestamp 1626908933
transform 1 0 9312 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_46
timestamp 1626908933
transform 1 0 8928 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_166
timestamp 1626908933
transform 1 0 8928 0 -1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_864
timestamp 1626908933
transform 1 0 9936 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_362
timestamp 1626908933
transform 1 0 9936 0 1 5661
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_136
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_17
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_136
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_17
timestamp 1626908933
transform 1 0 10100 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_63
timestamp 1626908933
transform -1 0 11424 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_62
timestamp 1626908933
transform -1 0 10752 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_29
timestamp 1626908933
transform -1 0 11424 0 -1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_28
timestamp 1626908933
transform -1 0 10752 0 -1 6660
box -38 -49 710 715
use L1M1_PR  L1M1_PR_858
timestamp 1626908933
transform 1 0 11472 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_356
timestamp 1626908933
transform 1 0 11472 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_766
timestamp 1626908933
transform 1 0 11472 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_301
timestamp 1626908933
transform 1 0 11472 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_227
timestamp 1626908933
transform 1 0 11616 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_57
timestamp 1626908933
transform 1 0 11616 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_135
timestamp 1626908933
transform 1 0 11424 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_22
timestamp 1626908933
transform 1 0 11424 0 -1 6660
box -38 -49 230 715
use L1M1_PR  L1M1_PR_785
timestamp 1626908933
transform 1 0 11856 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_283
timestamp 1626908933
transform 1 0 11856 0 1 5661
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_119
timestamp 1626908933
transform 1 0 11712 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_16
timestamp 1626908933
transform 1 0 11712 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_45
timestamp 1626908933
transform 1 0 12480 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_127
timestamp 1626908933
transform 1 0 12480 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_232
timestamp 1626908933
transform 1 0 12336 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_697
timestamp 1626908933
transform 1 0 12336 0 1 5661
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_6
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_125
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_6
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_125
timestamp 1626908933
transform 1 0 12500 0 1 5994
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_21
timestamp 1626908933
transform 1 0 12576 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_134
timestamp 1626908933
transform 1 0 12576 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_56
timestamp 1626908933
transform 1 0 12768 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_226
timestamp 1626908933
transform 1 0 12768 0 -1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_372
timestamp 1626908933
transform 1 0 12816 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_837
timestamp 1626908933
transform 1 0 12816 0 1 5883
box -32 -32 32 32
use M2M3_PR  M2M3_PR_21
timestamp 1626908933
transform 1 0 12816 0 1 5893
box -33 -37 33 37
use M2M3_PR  M2M3_PR_63
timestamp 1626908933
transform 1 0 12816 0 1 5893
box -33 -37 33 37
use L1M1_PR  L1M1_PR_391
timestamp 1626908933
transform 1 0 13200 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_893
timestamp 1626908933
transform 1 0 13200 0 1 5883
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_9
timestamp 1626908933
transform 1 0 13632 0 -1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_38
timestamp 1626908933
transform 1 0 13632 0 -1 6660
box -38 -49 326 715
use M1M2_PR  M1M2_PR_335
timestamp 1626908933
transform 1 0 13584 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_375
timestamp 1626908933
transform 1 0 13584 0 1 5439
box -32 -32 32 32
use M1M2_PR  M1M2_PR_800
timestamp 1626908933
transform 1 0 13584 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_840
timestamp 1626908933
transform 1 0 13584 0 1 5439
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_6
timestamp 1626908933
transform 1 0 12864 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_109
timestamp 1626908933
transform 1 0 12864 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_290
timestamp 1626908933
transform 1 0 13920 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_120
timestamp 1626908933
transform 1 0 13920 0 -1 6660
box -38 -49 134 715
use M2M3_PR  M2M3_PR_74
timestamp 1626908933
transform 1 0 240 0 1 6747
box -33 -37 33 37
use M2M3_PR  M2M3_PR_73
timestamp 1626908933
transform 1 0 240 0 1 6259
box -33 -37 33 37
use M2M3_PR  M2M3_PR_32
timestamp 1626908933
transform 1 0 240 0 1 6747
box -33 -37 33 37
use M2M3_PR  M2M3_PR_31
timestamp 1626908933
transform 1 0 240 0 1 6259
box -33 -37 33 37
use M1M2_PR  M1M2_PR_847
timestamp 1626908933
transform 1 0 240 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_382
timestamp 1626908933
transform 1 0 240 0 1 6105
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_291
timestamp 1626908933
transform 1 0 192 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_121
timestamp 1626908933
transform 1 0 192 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_126
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_44
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_184
timestamp 1626908933
transform 1 0 0 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_71
timestamp 1626908933
transform 1 0 0 0 1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_6
timestamp 1626908933
transform 1 0 912 0 1 6179
box -32 -32 32 32
use M1M2_PR  M1M2_PR_471
timestamp 1626908933
transform 1 0 912 0 1 6179
box -32 -32 32 32
use L1M1_PR  L1M1_PR_5
timestamp 1626908933
transform 1 0 912 0 1 6179
box -29 -23 29 23
use L1M1_PR  L1M1_PR_507
timestamp 1626908933
transform 1 0 912 0 1 6179
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_88
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_191
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_430
timestamp 1626908933
transform 1 0 1488 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_932
timestamp 1626908933
transform 1 0 1488 0 1 6105
box -29 -23 29 23
use M1M2_PR  M1M2_PR_340
timestamp 1626908933
transform 1 0 1104 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_805
timestamp 1626908933
transform 1 0 1104 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_172
timestamp 1626908933
transform 1 0 1104 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_674
timestamp 1626908933
transform 1 0 1104 0 1 6253
box -29 -23 29 23
use M1M2_PR  M1M2_PR_216
timestamp 1626908933
transform 1 0 1296 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_681
timestamp 1626908933
transform 1 0 1296 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_11
timestamp 1626908933
transform 1 0 1776 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_476
timestamp 1626908933
transform 1 0 1776 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_10
timestamp 1626908933
transform 1 0 1680 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_512
timestamp 1626908933
transform 1 0 1680 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_212
timestamp 1626908933
transform 1 0 1872 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_677
timestamp 1626908933
transform 1 0 1872 0 1 6401
box -32 -32 32 32
use L1M1_PR  L1M1_PR_263
timestamp 1626908933
transform 1 0 1872 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_493
timestamp 1626908933
transform 1 0 1968 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_765
timestamp 1626908933
transform 1 0 1872 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_995
timestamp 1626908933
transform 1 0 1968 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_396
timestamp 1626908933
transform 1 0 1200 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_898
timestamp 1626908933
transform 1 0 1200 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_15
timestamp 1626908933
transform 1 0 1488 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_480
timestamp 1626908933
transform 1 0 1488 0 1 6549
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_114
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_233
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_114
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_233
timestamp 1626908933
transform 1 0 1700 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_66
timestamp 1626908933
transform -1 0 3072 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_29
timestamp 1626908933
transform -1 0 3072 0 1 6660
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_887
timestamp 1626908933
transform 1 0 2832 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_847
timestamp 1626908933
transform 1 0 2256 0 1 6475
box -29 -23 29 23
use L1M1_PR  L1M1_PR_385
timestamp 1626908933
transform 1 0 2832 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_345
timestamp 1626908933
transform 1 0 2256 0 1 6475
box -29 -23 29 23
use M1M2_PR  M1M2_PR_919
timestamp 1626908933
transform 1 0 2064 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_619
timestamp 1626908933
transform 1 0 2736 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_454
timestamp 1626908933
transform 1 0 2064 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_154
timestamp 1626908933
transform 1 0 2736 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_846
timestamp 1626908933
transform 1 0 3216 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_344
timestamp 1626908933
transform 1 0 3216 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_790
timestamp 1626908933
transform 1 0 3504 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_325
timestamp 1626908933
transform 1 0 3504 0 1 6327
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_225
timestamp 1626908933
transform 1 0 3072 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_55
timestamp 1626908933
transform 1 0 3072 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_169
timestamp 1626908933
transform 1 0 3168 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_66
timestamp 1626908933
transform 1 0 3168 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_224
timestamp 1626908933
transform 1 0 3936 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_54
timestamp 1626908933
transform 1 0 3936 0 1 6660
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_223
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_104
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_223
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_104
timestamp 1626908933
transform 1 0 4100 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_292
timestamp 1626908933
transform 1 0 4032 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_122
timestamp 1626908933
transform 1 0 4032 0 1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_634
timestamp 1626908933
transform 1 0 4368 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_513
timestamp 1626908933
transform 1 0 4368 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_132
timestamp 1626908933
transform 1 0 4368 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_11
timestamp 1626908933
transform 1 0 4368 0 1 6549
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_223
timestamp 1626908933
transform 1 0 4416 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_53
timestamp 1626908933
transform 1 0 4416 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_32
timestamp 1626908933
transform 1 0 4128 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_3
timestamp 1626908933
transform 1 0 4128 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_72
timestamp 1626908933
transform 1 0 4512 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_192
timestamp 1626908933
transform 1 0 4512 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_43
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_125
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_52
timestamp 1626908933
transform 1 0 4896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_222
timestamp 1626908933
transform 1 0 4896 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_85
timestamp 1626908933
transform 1 0 5616 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_126
timestamp 1626908933
transform 1 0 5424 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_127
timestamp 1626908933
transform 1 0 5424 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_550
timestamp 1626908933
transform 1 0 5616 0 1 6845
box -32 -32 32 32
use M1M2_PR  M1M2_PR_591
timestamp 1626908933
transform 1 0 5424 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_592
timestamp 1626908933
transform 1 0 5424 0 1 6327
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_52
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_155
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_34
timestamp 1626908933
transform -1 0 6528 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_0
timestamp 1626908933
transform -1 0 6528 0 1 6660
box -38 -49 710 715
use L1M1_PR  L1M1_PR_636
timestamp 1626908933
transform 1 0 5808 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_633
timestamp 1626908933
transform 1 0 5808 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_134
timestamp 1626908933
transform 1 0 5808 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_131
timestamp 1626908933
transform 1 0 5808 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_128
timestamp 1626908933
transform 1 0 6288 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_593
timestamp 1626908933
transform 1 0 6288 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_130
timestamp 1626908933
transform 1 0 6096 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_632
timestamp 1626908933
transform 1 0 6096 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_686
timestamp 1626908933
transform 1 0 6384 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_684
timestamp 1626908933
transform 1 0 6480 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_184
timestamp 1626908933
transform 1 0 6384 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_182
timestamp 1626908933
transform 1 0 6480 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_626
timestamp 1626908933
transform 1 0 6384 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_624
timestamp 1626908933
transform 1 0 6672 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_161
timestamp 1626908933
transform 1 0 6384 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_159
timestamp 1626908933
transform 1 0 6672 0 1 6327
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_213
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_94
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_213
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_94
timestamp 1626908933
transform 1 0 6500 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_185
timestamp 1626908933
transform 1 0 6528 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_72
timestamp 1626908933
transform 1 0 6528 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_4
timestamp 1626908933
transform 1 0 6720 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_38
timestamp 1626908933
transform 1 0 6720 0 1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_125
timestamp 1626908933
transform 1 0 6960 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_590
timestamp 1626908933
transform 1 0 6960 0 1 6549
box -32 -32 32 32
use L1M1_PR  L1M1_PR_179
timestamp 1626908933
transform 1 0 7056 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_180
timestamp 1626908933
transform 1 0 6768 0 1 6475
box -29 -23 29 23
use L1M1_PR  L1M1_PR_681
timestamp 1626908933
transform 1 0 7056 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_682
timestamp 1626908933
transform 1 0 6768 0 1 6475
box -29 -23 29 23
use L1M1_PR  L1M1_PR_680
timestamp 1626908933
transform 1 0 7152 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_178
timestamp 1626908933
transform 1 0 7152 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_638
timestamp 1626908933
transform 1 0 7440 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_136
timestamp 1626908933
transform 1 0 7440 0 1 6549
box -29 -23 29 23
use M1M2_PR  M1M2_PR_622
timestamp 1626908933
transform 1 0 7344 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_621
timestamp 1626908933
transform 1 0 7344 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_157
timestamp 1626908933
transform 1 0 7344 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_156
timestamp 1626908933
transform 1 0 7344 0 1 6771
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_293
timestamp 1626908933
transform 1 0 7392 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_123
timestamp 1626908933
transform 1 0 7392 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_6
timestamp 1626908933
transform -1 0 8160 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_40
timestamp 1626908933
transform -1 0 8160 0 1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_596
timestamp 1626908933
transform 1 0 7728 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_131
timestamp 1626908933
transform 1 0 7728 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_55
timestamp 1626908933
transform -1 0 8832 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_21
timestamp 1626908933
transform -1 0 8832 0 1 6660
box -38 -49 710 715
use L1M1_PR  L1M1_PR_679
timestamp 1626908933
transform 1 0 8208 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_177
timestamp 1626908933
transform 1 0 8208 0 1 6771
box -29 -23 29 23
use M1M2_PR  M1M2_PR_523
timestamp 1626908933
transform 1 0 8400 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_58
timestamp 1626908933
transform 1 0 8400 0 1 6105
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_203
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_84
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_203
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_84
timestamp 1626908933
transform 1 0 8900 0 1 6660
box -100 -49 100 49
use L1M1_PR  L1M1_PR_584
timestamp 1626908933
transform 1 0 8976 0 1 6845
box -29 -23 29 23
use L1M1_PR  L1M1_PR_82
timestamp 1626908933
transform 1 0 8976 0 1 6845
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_186
timestamp 1626908933
transform 1 0 8832 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_73
timestamp 1626908933
transform 1 0 8832 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_55
timestamp 1626908933
transform 1 0 9024 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_26
timestamp 1626908933
transform 1 0 9024 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_30
timestamp 1626908933
transform 1 0 9312 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_64
timestamp 1626908933
transform 1 0 9312 0 1 6660
box -38 -49 710 715
use L1M1_PR  L1M1_PR_724
timestamp 1626908933
transform 1 0 9936 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_222
timestamp 1626908933
transform 1 0 9936 0 1 6771
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_124
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_42
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_178
timestamp 1626908933
transform 1 0 10128 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_179
timestamp 1626908933
transform 1 0 10128 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_643
timestamp 1626908933
transform 1 0 10128 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_644
timestamp 1626908933
transform 1 0 10128 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_220
timestamp 1626908933
transform 1 0 10128 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_221
timestamp 1626908933
transform 1 0 10416 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_722
timestamp 1626908933
transform 1 0 10128 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_723
timestamp 1626908933
transform 1 0 10416 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_726
timestamp 1626908933
transform 1 0 10512 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_224
timestamp 1626908933
transform 1 0 10512 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_642
timestamp 1626908933
transform 1 0 10512 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_521
timestamp 1626908933
transform 1 0 10512 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_177
timestamp 1626908933
transform 1 0 10512 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_56
timestamp 1626908933
transform 1 0 10512 0 1 6105
box -32 -32 32 32
use L1M1_PR  L1M1_PR_725
timestamp 1626908933
transform 1 0 10800 0 1 6475
box -29 -23 29 23
use L1M1_PR  L1M1_PR_223
timestamp 1626908933
transform 1 0 10800 0 1 6475
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_221
timestamp 1626908933
transform 1 0 10752 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_51
timestamp 1626908933
transform 1 0 10752 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_147
timestamp 1626908933
transform 1 0 10848 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_27
timestamp 1626908933
transform 1 0 10848 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_27
timestamp 1626908933
transform -1 0 10752 0 1 6660
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_61
timestamp 1626908933
transform -1 0 10752 0 1 6660
box -38 -49 710 715
use M1M2_PR  M1M2_PR_183
timestamp 1626908933
transform 1 0 10992 0 1 6253
box -32 -32 32 32
use M1M2_PR  M1M2_PR_648
timestamp 1626908933
transform 1 0 10992 0 1 6253
box -32 -32 32 32
use L1M1_PR  L1M1_PR_226
timestamp 1626908933
transform 1 0 11088 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_228
timestamp 1626908933
transform 1 0 11088 0 1 6253
box -29 -23 29 23
use L1M1_PR  L1M1_PR_728
timestamp 1626908933
transform 1 0 11088 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_730
timestamp 1626908933
transform 1 0 11088 0 1 6253
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_50
timestamp 1626908933
transform 1 0 11232 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_220
timestamp 1626908933
transform 1 0 11232 0 1 6660
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_74
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_193
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_74
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_193
timestamp 1626908933
transform 1 0 11300 0 1 6660
box -100 -49 100 49
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_56
timestamp 1626908933
transform 1 0 11328 0 1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_19
timestamp 1626908933
transform 1 0 11328 0 1 6660
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_645
timestamp 1626908933
transform 1 0 12048 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_180
timestamp 1626908933
transform 1 0 12048 0 1 6327
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_122
timestamp 1626908933
transform 1 0 13248 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_2
timestamp 1626908933
transform 1 0 13248 0 1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_56
timestamp 1626908933
transform 1 0 13584 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_558
timestamp 1626908933
transform 1 0 13584 0 1 6105
box -29 -23 29 23
use M2M3_PR  M2M3_PR_4
timestamp 1626908933
transform 1 0 13584 0 1 6503
box -33 -37 33 37
use M2M3_PR  M2M3_PR_46
timestamp 1626908933
transform 1 0 13584 0 1 6503
box -33 -37 33 37
use L1M1_PR  L1M1_PR_667
timestamp 1626908933
transform 1 0 13776 0 1 6105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_165
timestamp 1626908933
transform 1 0 13776 0 1 6105
box -29 -23 29 23
use M1M2_PR  M1M2_PR_617
timestamp 1626908933
transform 1 0 13776 0 1 6105
box -32 -32 32 32
use M1M2_PR  M1M2_PR_152
timestamp 1626908933
transform 1 0 13776 0 1 6105
box -32 -32 32 32
use prbs_generator_syn_VIA10  prbs_generator_syn_VIA10_1
timestamp 1626908933
transform 1 0 13700 0 1 6681
box -100 -28 100 28
use prbs_generator_syn_VIA10  prbs_generator_syn_VIA10_0
timestamp 1626908933
transform 1 0 13700 0 1 6681
box -100 -28 100 28
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_12
timestamp 1626908933
transform 1 0 13700 0 1 6676
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_4
timestamp 1626908933
transform 1 0 13700 0 1 6676
box -100 -33 100 33
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_123
timestamp 1626908933
transform 1 0 13632 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_41
timestamp 1626908933
transform 1 0 13632 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_74
timestamp 1626908933
transform 1 0 13728 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_187
timestamp 1626908933
transform 1 0 13728 0 1 6660
box -38 -49 230 715
use L1M1_PR  L1M1_PR_915
timestamp 1626908933
transform 1 0 13872 0 1 6401
box -29 -23 29 23
use L1M1_PR  L1M1_PR_413
timestamp 1626908933
transform 1 0 13872 0 1 6401
box -29 -23 29 23
use M1M2_PR  M1M2_PR_824
timestamp 1626908933
transform 1 0 13872 0 1 6401
box -32 -32 32 32
use M1M2_PR  M1M2_PR_359
timestamp 1626908933
transform 1 0 13872 0 1 6401
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_294
timestamp 1626908933
transform 1 0 13920 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_124
timestamp 1626908933
transform 1 0 13920 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_49
timestamp 1626908933
transform 1 0 0 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_219
timestamp 1626908933
transform 1 0 0 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_339
timestamp 1626908933
transform 1 0 144 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_383
timestamp 1626908933
transform 1 0 48 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_804
timestamp 1626908933
transform 1 0 144 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_848
timestamp 1626908933
transform 1 0 48 0 1 7437
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_60
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_179
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_60
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_179
timestamp 1626908933
transform 1 0 500 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_97
timestamp 1626908933
transform 1 0 96 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_200
timestamp 1626908933
transform 1 0 96 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_48
timestamp 1626908933
transform 1 0 1248 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_218
timestamp 1626908933
transform 1 0 1248 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_18
timestamp 1626908933
transform 1 0 912 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_483
timestamp 1626908933
transform 1 0 912 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_16
timestamp 1626908933
transform 1 0 1296 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_431
timestamp 1626908933
transform 1 0 1296 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_518
timestamp 1626908933
transform 1 0 1296 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_933
timestamp 1626908933
transform 1 0 1296 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_108
timestamp 1626908933
transform 1 0 864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_228
timestamp 1626908933
transform 1 0 864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_27
timestamp 1626908933
transform 1 0 1344 0 -1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_59
timestamp 1626908933
transform 1 0 1344 0 -1 7992
box -38 -49 710 715
use L1M1_PR  L1M1_PR_845
timestamp 1626908933
transform 1 0 1968 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_343
timestamp 1626908933
transform 1 0 1968 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_40
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_122
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_92
timestamp 1626908933
transform 1 0 2112 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_212
timestamp 1626908933
transform 1 0 2112 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_47
timestamp 1626908933
transform 1 0 2016 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_217
timestamp 1626908933
transform 1 0 2016 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_844
timestamp 1626908933
transform 1 0 2640 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_342
timestamp 1626908933
transform 1 0 2640 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_752
timestamp 1626908933
transform 1 0 2544 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_287
timestamp 1626908933
transform 1 0 2544 0 1 6993
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_168
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_49
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_168
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_49
timestamp 1626908933
transform 1 0 2900 0 1 7326
box -100 -49 100 49
use M1M2_PR  M1M2_PR_751
timestamp 1626908933
transform 1 0 2544 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_286
timestamp 1626908933
transform 1 0 2544 0 1 7437
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_69
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_172
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_885
timestamp 1626908933
transform 1 0 3024 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_383
timestamp 1626908933
transform 1 0 3024 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_789
timestamp 1626908933
transform 1 0 3504 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_467
timestamp 1626908933
transform 1 0 3888 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_324
timestamp 1626908933
transform 1 0 3504 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2
timestamp 1626908933
transform 1 0 3888 0 1 6919
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_188
timestamp 1626908933
transform 1 0 3360 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_75
timestamp 1626908933
transform 1 0 3360 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_65
timestamp 1626908933
transform 1 0 3552 0 -1 7992
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_28
timestamp 1626908933
transform 1 0 3552 0 -1 7992
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_897
timestamp 1626908933
transform 1 0 4464 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_504
timestamp 1626908933
transform 1 0 4176 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_395
timestamp 1626908933
transform 1 0 4464 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2
timestamp 1626908933
transform 1 0 4176 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_112
timestamp 1626908933
transform 1 0 4944 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_577
timestamp 1626908933
transform 1 0 4944 0 1 6919
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_38
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_157
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_38
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_157
timestamp 1626908933
transform 1 0 5300 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_46
timestamp 1626908933
transform 1 0 5472 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_216
timestamp 1626908933
transform 1 0 5472 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_51
timestamp 1626908933
transform 1 0 5568 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_154
timestamp 1626908933
transform 1 0 5568 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_611
timestamp 1626908933
transform 1 0 5808 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_109
timestamp 1626908933
transform 1 0 5808 0 1 6919
box -29 -23 29 23
use M1M2_PR  M1M2_PR_115
timestamp 1626908933
transform 1 0 6000 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_580
timestamp 1626908933
transform 1 0 6000 0 1 7067
box -32 -32 32 32
use L1M1_PR  L1M1_PR_112
timestamp 1626908933
transform 1 0 6192 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_113
timestamp 1626908933
transform 1 0 6192 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_614
timestamp 1626908933
transform 1 0 6192 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_615
timestamp 1626908933
transform 1 0 6192 0 1 7067
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_42
timestamp 1626908933
transform 1 0 6720 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_145
timestamp 1626908933
transform 1 0 6720 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_62
timestamp 1626908933
transform 1 0 6336 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_182
timestamp 1626908933
transform 1 0 6336 0 -1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_124
timestamp 1626908933
transform 1 0 6960 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_589
timestamp 1626908933
transform 1 0 6960 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_128
timestamp 1626908933
transform 1 0 7056 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_129
timestamp 1626908933
transform 1 0 6960 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_630
timestamp 1626908933
transform 1 0 7056 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_631
timestamp 1626908933
transform 1 0 6960 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_123
timestamp 1626908933
transform 1 0 7248 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_588
timestamp 1626908933
transform 1 0 7248 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_126
timestamp 1626908933
transform 1 0 7152 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_628
timestamp 1626908933
transform 1 0 7152 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_629
timestamp 1626908933
transform 1 0 7440 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_127
timestamp 1626908933
transform 1 0 7440 0 1 6993
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_146
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_27
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_146
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_27
timestamp 1626908933
transform 1 0 7700 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_133
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_20
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_121
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_39
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_45
timestamp 1626908933
transform 1 0 7776 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_215
timestamp 1626908933
transform 1 0 7776 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_130
timestamp 1626908933
transform 1 0 7728 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_595
timestamp 1626908933
transform 1 0 7728 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_135
timestamp 1626908933
transform 1 0 7824 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_138
timestamp 1626908933
transform 1 0 7920 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_637
timestamp 1626908933
transform 1 0 7824 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_640
timestamp 1626908933
transform 1 0 7920 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_34
timestamp 1626908933
transform 1 0 7872 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_137
timestamp 1626908933
transform 1 0 7872 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_698
timestamp 1626908933
transform 1 0 8592 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_696
timestamp 1626908933
transform 1 0 8496 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_196
timestamp 1626908933
transform 1 0 8592 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_194
timestamp 1626908933
transform 1 0 8496 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_630
timestamp 1626908933
transform 1 0 8592 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_598
timestamp 1626908933
transform 1 0 8400 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_165
timestamp 1626908933
transform 1 0 8592 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_133
timestamp 1626908933
transform 1 0 8400 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_629
timestamp 1626908933
transform 1 0 8592 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_164
timestamp 1626908933
transform 1 0 8592 0 1 7437
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_47
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_18
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_195
timestamp 1626908933
transform 1 0 8784 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_697
timestamp 1626908933
transform 1 0 8784 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_162
timestamp 1626908933
transform 1 0 8880 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_163
timestamp 1626908933
transform 1 0 8880 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_627
timestamp 1626908933
transform 1 0 8880 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_628
timestamp 1626908933
transform 1 0 8880 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_230
timestamp 1626908933
transform 1 0 9168 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_419
timestamp 1626908933
transform 1 0 8976 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_732
timestamp 1626908933
transform 1 0 9168 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_921
timestamp 1626908933
transform 1 0 8976 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_923
timestamp 1626908933
transform 1 0 9264 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_421
timestamp 1626908933
transform 1 0 9264 0 1 6919
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_295
timestamp 1626908933
transform 1 0 9312 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_125
timestamp 1626908933
transform 1 0 9312 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_734
timestamp 1626908933
transform 1 0 9648 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_731
timestamp 1626908933
transform 1 0 9648 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_695
timestamp 1626908933
transform 1 0 9552 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_232
timestamp 1626908933
transform 1 0 9648 0 1 7067
box -29 -23 29 23
use L1M1_PR  L1M1_PR_229
timestamp 1626908933
transform 1 0 9648 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_193
timestamp 1626908933
transform 1 0 9552 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_650
timestamp 1626908933
transform 1 0 9552 0 1 7067
box -32 -32 32 32
use M1M2_PR  M1M2_PR_185
timestamp 1626908933
transform 1 0 9552 0 1 7067
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_48
timestamp 1626908933
transform 1 0 9408 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_19
timestamp 1626908933
transform 1 0 9408 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_3
timestamp 1626908933
transform 1 0 8928 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_10
timestamp 1626908933
transform 1 0 8928 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_214
timestamp 1626908933
transform 1 0 9696 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_44
timestamp 1626908933
transform 1 0 9696 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_129
timestamp 1626908933
transform 1 0 9792 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_26
timestamp 1626908933
transform 1 0 9792 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_111
timestamp 1626908933
transform 1 0 10320 0 1 7141
box -29 -23 29 23
use L1M1_PR  L1M1_PR_613
timestamp 1626908933
transform 1 0 10320 0 1 7141
box -29 -23 29 23
use M1M2_PR  M1M2_PR_175
timestamp 1626908933
transform 1 0 10416 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_640
timestamp 1626908933
transform 1 0 10416 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_218
timestamp 1626908933
transform 1 0 10416 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_720
timestamp 1626908933
transform 1 0 10416 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_176
timestamp 1626908933
transform 1 0 10512 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_641
timestamp 1626908933
transform 1 0 10512 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_219
timestamp 1626908933
transform 1 0 10512 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_721
timestamp 1626908933
transform 1 0 10512 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_357
timestamp 1626908933
transform 1 0 11376 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_859
timestamp 1626908933
transform 1 0 11376 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_300
timestamp 1626908933
transform 1 0 11664 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_765
timestamp 1626908933
transform 1 0 11664 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_323
timestamp 1626908933
transform 1 0 11760 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_825
timestamp 1626908933
transform 1 0 11760 0 1 6993
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_16
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_135
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_16
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_135
timestamp 1626908933
transform 1 0 10100 0 1 7326
box -100 -49 100 49
use M1M2_PR  M1M2_PR_54
timestamp 1626908933
transform 1 0 10704 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_174
timestamp 1626908933
transform 1 0 10608 0 1 7511
box -32 -32 32 32
use M1M2_PR  M1M2_PR_519
timestamp 1626908933
transform 1 0 10704 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_639
timestamp 1626908933
transform 1 0 10608 0 1 7511
box -32 -32 32 32
use L1M1_PR  L1M1_PR_54
timestamp 1626908933
transform 1 0 10704 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_556
timestamp 1626908933
transform 1 0 10704 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_54
timestamp 1626908933
transform -1 0 12480 0 -1 7992
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_17
timestamp 1626908933
transform -1 0 12480 0 -1 7992
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_269
timestamp 1626908933
transform 1 0 12144 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_734
timestamp 1626908933
transform 1 0 12144 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_38
timestamp 1626908933
transform 1 0 12480 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_120
timestamp 1626908933
transform 1 0 12480 0 -1 7992
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_5
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_124
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_5
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_124
timestamp 1626908933
transform 1 0 12500 0 1 7326
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_5
timestamp 1626908933
transform 1 0 12576 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_108
timestamp 1626908933
transform 1 0 12576 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_44
timestamp 1626908933
transform 1 0 13488 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_371
timestamp 1626908933
transform 1 0 13392 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_509
timestamp 1626908933
transform 1 0 13488 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_836
timestamp 1626908933
transform 1 0 13392 0 1 6919
box -32 -32 32 32
use L1M1_PR  L1M1_PR_46
timestamp 1626908933
transform 1 0 13104 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_548
timestamp 1626908933
transform 1 0 13104 0 1 7215
box -29 -23 29 23
use M2M3_PR  M2M3_PR_20
timestamp 1626908933
transform 1 0 13392 0 1 7113
box -33 -37 33 37
use M2M3_PR  M2M3_PR_62
timestamp 1626908933
transform 1 0 13392 0 1 7113
box -33 -37 33 37
use M1M2_PR  M1M2_PR_369
timestamp 1626908933
transform 1 0 13104 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_834
timestamp 1626908933
transform 1 0 13104 0 1 7585
box -32 -32 32 32
use L1M1_PR  L1M1_PR_217
timestamp 1626908933
transform 1 0 13584 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_719
timestamp 1626908933
transform 1 0 13584 0 1 7437
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_31
timestamp 1626908933
transform -1 0 14016 0 -1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_65
timestamp 1626908933
transform -1 0 14016 0 -1 7992
box -38 -49 710 715
use L1M1_PR  L1M1_PR_738
timestamp 1626908933
transform 1 0 13680 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_236
timestamp 1626908933
transform 1 0 13680 0 1 7585
box -29 -23 29 23
use M1M2_PR  M1M2_PR_653
timestamp 1626908933
transform 1 0 13968 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_188
timestamp 1626908933
transform 1 0 13968 0 1 7585
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_296
timestamp 1626908933
transform 1 0 192 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_126
timestamp 1626908933
transform 1 0 192 0 1 7992
box -38 -49 134 715
use M2M3_PR  M2M3_PR_75
timestamp 1626908933
transform 1 0 240 0 1 8211
box -33 -37 33 37
use M2M3_PR  M2M3_PR_33
timestamp 1626908933
transform 1 0 240 0 1 8211
box -33 -37 33 37
use M1M2_PR  M1M2_PR_850
timestamp 1626908933
transform 1 0 240 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_849
timestamp 1626908933
transform 1 0 336 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_385
timestamp 1626908933
transform 1 0 240 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_384
timestamp 1626908933
transform 1 0 336 0 1 8103
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_119
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_37
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_189
timestamp 1626908933
transform 1 0 0 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_132
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_76
timestamp 1626908933
transform 1 0 0 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_19
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_87
timestamp 1626908933
transform 1 0 576 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_190
timestamp 1626908933
transform 1 0 576 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_515
timestamp 1626908933
transform 1 0 1488 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_13
timestamp 1626908933
transform 1 0 1488 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_479
timestamp 1626908933
transform 1 0 1488 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_14
timestamp 1626908933
transform 1 0 1488 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_767
timestamp 1626908933
transform 1 0 1680 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_265
timestamp 1626908933
transform 1 0 1680 0 1 7659
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_232
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_113
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_232
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_113
timestamp 1626908933
transform 1 0 1700 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_934
timestamp 1626908933
transform 1 0 1392 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_432
timestamp 1626908933
transform 1 0 1392 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_482
timestamp 1626908933
transform 1 0 912 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_17
timestamp 1626908933
transform 1 0 912 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_517
timestamp 1626908933
transform 1 0 1392 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_15
timestamp 1626908933
transform 1 0 1392 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_766
timestamp 1626908933
transform 1 0 1680 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_264
timestamp 1626908933
transform 1 0 1680 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_680
timestamp 1626908933
transform 1 0 1680 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_215
timestamp 1626908933
transform 1 0 1680 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_26
timestamp 1626908933
transform 1 0 1344 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_58
timestamp 1626908933
transform 1 0 1344 0 1 7992
box -38 -49 710 715
use L1M1_PR  L1M1_PR_998
timestamp 1626908933
transform 1 0 1776 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_997
timestamp 1626908933
transform 1 0 1776 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_843
timestamp 1626908933
transform 1 0 1968 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_496
timestamp 1626908933
transform 1 0 1776 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_495
timestamp 1626908933
transform 1 0 1776 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_341
timestamp 1626908933
transform 1 0 1968 0 1 8177
box -29 -23 29 23
use M1M2_PR  M1M2_PR_676
timestamp 1626908933
transform 1 0 1872 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_211
timestamp 1626908933
transform 1 0 1872 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_22
timestamp 1626908933
transform 1 0 2640 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_453
timestamp 1626908933
transform 1 0 2064 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_487
timestamp 1626908933
transform 1 0 2640 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_918
timestamp 1626908933
transform 1 0 2064 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_935
timestamp 1626908933
transform 1 0 2448 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_433
timestamp 1626908933
transform 1 0 2448 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_917
timestamp 1626908933
transform 1 0 2064 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_452
timestamp 1626908933
transform 1 0 2064 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_521
timestamp 1626908933
transform 1 0 2544 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_19
timestamp 1626908933
transform 1 0 2544 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_763
timestamp 1626908933
transform 1 0 2736 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_261
timestamp 1626908933
transform 1 0 2736 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_672
timestamp 1626908933
transform 1 0 2736 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_486
timestamp 1626908933
transform 1 0 2640 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_207
timestamp 1626908933
transform 1 0 2736 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_21
timestamp 1626908933
transform 1 0 2640 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_994
timestamp 1626908933
transform 1 0 2832 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_492
timestamp 1626908933
transform 1 0 2832 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_91
timestamp 1626908933
transform 1 0 2016 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_211
timestamp 1626908933
transform 1 0 2016 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_25
timestamp 1626908933
transform 1 0 2400 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_57
timestamp 1626908933
transform 1 0 2400 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_43
timestamp 1626908933
transform 1 0 3072 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_213
timestamp 1626908933
transform 1 0 3072 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_284
timestamp 1626908933
transform 1 0 3312 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_285
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_323
timestamp 1626908933
transform 1 0 3600 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_749
timestamp 1626908933
transform 1 0 3312 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_750
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_788
timestamp 1626908933
transform 1 0 3600 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_381
timestamp 1626908933
transform 1 0 3600 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_883
timestamp 1626908933
transform 1 0 3600 0 1 7659
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_65
timestamp 1626908933
transform 1 0 3168 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_168
timestamp 1626908933
transform 1 0 3168 0 1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_842
timestamp 1626908933
transform 1 0 3984 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_340
timestamp 1626908933
transform 1 0 3984 0 1 7733
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_131
timestamp 1626908933
transform 1 0 3936 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_18
timestamp 1626908933
transform 1 0 3936 0 1 7992
box -38 -49 230 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_222
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_103
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_222
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_103
timestamp 1626908933
transform 1 0 4100 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_212
timestamp 1626908933
transform 1 0 4128 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_42
timestamp 1626908933
transform 1 0 4128 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_161
timestamp 1626908933
transform 1 0 4224 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_58
timestamp 1626908933
transform 1 0 4224 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_36
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_118
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_41
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_211
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_20
timestamp 1626908933
transform 1 0 5040 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_485
timestamp 1626908933
transform 1 0 5040 0 1 7881
box -32 -32 32 32
use L1M1_PR  L1M1_PR_17
timestamp 1626908933
transform 1 0 5136 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_519
timestamp 1626908933
transform 1 0 5136 0 1 7881
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_50
timestamp 1626908933
transform 1 0 5184 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_153
timestamp 1626908933
transform 1 0 5184 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_35
timestamp 1626908933
transform -1 0 6624 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_1
timestamp 1626908933
transform -1 0 6624 0 1 7992
box -38 -49 710 715
use M1M2_PR  M1M2_PR_114
timestamp 1626908933
transform 1 0 6000 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_579
timestamp 1626908933
transform 1 0 6000 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_114
timestamp 1626908933
transform 1 0 6000 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_116
timestamp 1626908933
transform 1 0 6288 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_616
timestamp 1626908933
transform 1 0 6000 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_618
timestamp 1626908933
transform 1 0 6288 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_127
timestamp 1626908933
transform 1 0 6624 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_297
timestamp 1626908933
transform 1 0 6624 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_115
timestamp 1626908933
transform 1 0 6672 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_617
timestamp 1626908933
transform 1 0 6672 0 1 8325
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_93
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_212
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_93
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_212
timestamp 1626908933
transform 1 0 6500 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_3
timestamp 1626908933
transform -1 0 7392 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_37
timestamp 1626908933
transform -1 0 7392 0 1 7992
box -38 -49 710 715
use M1M2_PR  M1M2_PR_121
timestamp 1626908933
transform 1 0 7056 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_122
timestamp 1626908933
transform 1 0 7248 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_586
timestamp 1626908933
transform 1 0 7056 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_587
timestamp 1626908933
transform 1 0 7248 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_124
timestamp 1626908933
transform 1 0 7056 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_125
timestamp 1626908933
transform 1 0 7152 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_626
timestamp 1626908933
transform 1 0 7056 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_627
timestamp 1626908933
transform 1 0 7152 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_77
timestamp 1626908933
transform 1 0 7392 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_190
timestamp 1626908933
transform 1 0 7392 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_41
timestamp 1626908933
transform 1 0 7584 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_7
timestamp 1626908933
transform 1 0 7584 0 1 7992
box -38 -49 710 715
use L1M1_PR  L1M1_PR_642
timestamp 1626908933
transform 1 0 7920 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_140
timestamp 1626908933
transform 1 0 7920 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_128
timestamp 1626908933
transform 1 0 8256 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_298
timestamp 1626908933
transform 1 0 8256 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_137
timestamp 1626908933
transform 1 0 8208 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_139
timestamp 1626908933
transform 1 0 8304 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_639
timestamp 1626908933
transform 1 0 8208 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_641
timestamp 1626908933
transform 1 0 8304 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_78
timestamp 1626908933
transform 1 0 8688 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_132
timestamp 1626908933
transform 1 0 8400 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_543
timestamp 1626908933
transform 1 0 8688 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_597
timestamp 1626908933
transform 1 0 8400 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_77
timestamp 1626908933
transform 1 0 8688 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_148
timestamp 1626908933
transform 1 0 8688 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_579
timestamp 1626908933
transform 1 0 8688 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_650
timestamp 1626908933
transform 1 0 8688 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_9
timestamp 1626908933
transform -1 0 9024 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_43
timestamp 1626908933
transform -1 0 9024 0 1 7992
box -38 -49 710 715
use M1M2_PR  M1M2_PR_74
timestamp 1626908933
transform 1 0 9456 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_539
timestamp 1626908933
transform 1 0 9456 0 1 7733
box -32 -32 32 32
use L1M1_PR  L1M1_PR_73
timestamp 1626908933
transform 1 0 9456 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_575
timestamp 1626908933
transform 1 0 9456 0 1 7733
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_83
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_202
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_83
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_202
timestamp 1626908933
transform 1 0 8900 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_147
timestamp 1626908933
transform 1 0 9072 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_174
timestamp 1626908933
transform 1 0 9360 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_176
timestamp 1626908933
transform 1 0 9456 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_649
timestamp 1626908933
transform 1 0 9072 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_676
timestamp 1626908933
transform 1 0 9360 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_678
timestamp 1626908933
transform 1 0 9456 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_16
timestamp 1626908933
transform -1 0 9696 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_50
timestamp 1626908933
transform -1 0 9696 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_78
timestamp 1626908933
transform 1 0 9696 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_191
timestamp 1626908933
transform 1 0 9696 0 1 7992
box -38 -49 230 715
use L1M1_PR  L1M1_PR_418
timestamp 1626908933
transform 1 0 9744 0 1 7881
box -29 -23 29 23
use L1M1_PR  L1M1_PR_920
timestamp 1626908933
transform 1 0 9744 0 1 7881
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_35
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_117
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_129
timestamp 1626908933
transform 1 0 9888 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_299
timestamp 1626908933
transform 1 0 9888 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_62
timestamp 1626908933
transform 1 0 9936 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_527
timestamp 1626908933
transform 1 0 9936 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_12
timestamp 1626908933
transform 1 0 10080 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_41
timestamp 1626908933
transform 1 0 10080 0 1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_63
timestamp 1626908933
transform 1 0 10128 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_175
timestamp 1626908933
transform 1 0 10224 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_565
timestamp 1626908933
transform 1 0 10128 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_677
timestamp 1626908933
transform 1 0 10224 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_555
timestamp 1626908933
transform 1 0 10704 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_53
timestamp 1626908933
transform 1 0 10704 0 1 8251
box -29 -23 29 23
use M1M2_PR  M1M2_PR_518
timestamp 1626908933
transform 1 0 10704 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_53
timestamp 1626908933
transform 1 0 10704 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_300
timestamp 1626908933
transform 1 0 10560 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_130
timestamp 1626908933
transform 1 0 10560 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_192
timestamp 1626908933
transform 1 0 10368 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_79
timestamp 1626908933
transform 1 0 10368 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_42
timestamp 1626908933
transform 1 0 10656 0 1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_13
timestamp 1626908933
transform 1 0 10656 0 1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_914
timestamp 1626908933
transform 1 0 10896 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_675
timestamp 1626908933
transform 1 0 10800 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_412
timestamp 1626908933
transform 1 0 10896 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_173
timestamp 1626908933
transform 1 0 10800 0 1 8177
box -29 -23 29 23
use M1M2_PR  M1M2_PR_823
timestamp 1626908933
transform 1 0 10896 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_657
timestamp 1626908933
transform 1 0 11088 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_358
timestamp 1626908933
transform 1 0 10896 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_192
timestamp 1626908933
transform 1 0 11088 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_193
timestamp 1626908933
transform 1 0 10944 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_80
timestamp 1626908933
transform 1 0 10944 0 1 7992
box -38 -49 230 715
use L1M1_PR  L1M1_PR_240
timestamp 1626908933
transform 1 0 11472 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_444
timestamp 1626908933
transform 1 0 11184 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_742
timestamp 1626908933
transform 1 0 11472 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_946
timestamp 1626908933
transform 1 0 11184 0 1 8103
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_73
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_192
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_73
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_192
timestamp 1626908933
transform 1 0 11300 0 1 7992
box -100 -49 100 49
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_14
timestamp 1626908933
transform 1 0 11136 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_46
timestamp 1626908933
transform 1 0 11136 0 1 7992
box -38 -49 710 715
use M1M2_PR  M1M2_PR_299
timestamp 1626908933
transform 1 0 11664 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_764
timestamp 1626908933
transform 1 0 11664 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_467
timestamp 1626908933
transform 1 0 11568 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_969
timestamp 1626908933
transform 1 0 11568 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_81
timestamp 1626908933
transform 1 0 11808 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_194
timestamp 1626908933
transform 1 0 11808 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_402
timestamp 1626908933
transform 1 0 11856 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_867
timestamp 1626908933
transform 1 0 11856 0 1 8177
box -32 -32 32 32
use L1M1_PR  L1M1_PR_317
timestamp 1626908933
transform 1 0 11760 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_819
timestamp 1626908933
transform 1 0 11760 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_265
timestamp 1626908933
transform 1 0 12048 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_730
timestamp 1626908933
transform 1 0 12048 0 1 7733
box -32 -32 32 32
use L1M1_PR  L1M1_PR_316
timestamp 1626908933
transform 1 0 12048 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_818
timestamp 1626908933
transform 1 0 12048 0 1 7733
box -29 -23 29 23
use M1M2_PR  M1M2_PR_264
timestamp 1626908933
transform 1 0 12048 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_268
timestamp 1626908933
transform 1 0 12144 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_729
timestamp 1626908933
transform 1 0 12048 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_733
timestamp 1626908933
transform 1 0 12144 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_322
timestamp 1626908933
transform 1 0 12144 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_824
timestamp 1626908933
transform 1 0 12144 0 1 8103
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_131
timestamp 1626908933
transform 1 0 12000 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_301
timestamp 1626908933
transform 1 0 12000 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_968
timestamp 1626908933
transform 1 0 12336 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_466
timestamp 1626908933
transform 1 0 12336 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_864
timestamp 1626908933
transform 1 0 12336 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_399
timestamp 1626908933
transform 1 0 12336 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_854
timestamp 1626908933
transform 1 0 12432 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_352
timestamp 1626908933
transform 1 0 12432 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_943
timestamp 1626908933
transform 1 0 12720 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_441
timestamp 1626908933
transform 1 0 12720 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_741
timestamp 1626908933
transform 1 0 12432 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_239
timestamp 1626908933
transform 1 0 12432 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_543
timestamp 1626908933
transform 1 0 12624 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_41
timestamp 1626908933
transform 1 0 12624 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_507
timestamp 1626908933
transform 1 0 12528 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_42
timestamp 1626908933
transform 1 0 12528 0 1 8325
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_17
timestamp 1626908933
transform -1 0 12768 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_49
timestamp 1626908933
transform -1 0 12768 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_82
timestamp 1626908933
transform 1 0 12768 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_195
timestamp 1626908933
transform 1 0 12768 0 1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_368
timestamp 1626908933
transform 1 0 13008 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_400
timestamp 1626908933
transform 1 0 12912 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_833
timestamp 1626908933
transform 1 0 13008 0 1 7881
box -32 -32 32 32
use M1M2_PR  M1M2_PR_865
timestamp 1626908933
transform 1 0 12912 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_46
timestamp 1626908933
transform 1 0 13392 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_511
timestamp 1626908933
transform 1 0 13392 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_237
timestamp 1626908933
transform 1 0 13296 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_462
timestamp 1626908933
transform 1 0 13200 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_739
timestamp 1626908933
transform 1 0 13296 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_964
timestamp 1626908933
transform 1 0 13200 0 1 8325
box -29 -23 29 23
use M2M3_PR  M2M3_PR_18
timestamp 1626908933
transform 1 0 13104 0 1 8333
box -33 -37 33 37
use M2M3_PR  M2M3_PR_60
timestamp 1626908933
transform 1 0 13104 0 1 8333
box -33 -37 33 37
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_16
timestamp 1626908933
transform -1 0 13632 0 1 7992
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_48
timestamp 1626908933
transform -1 0 13632 0 1 7992
box -38 -49 710 715
use M1M2_PR  M1M2_PR_187
timestamp 1626908933
transform 1 0 13488 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_652
timestamp 1626908933
transform 1 0 13488 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_234
timestamp 1626908933
transform 1 0 13680 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_736
timestamp 1626908933
transform 1 0 13680 0 1 7659
box -29 -23 29 23
use M2M3_PR  M2M3_PR_19
timestamp 1626908933
transform 1 0 13680 0 1 7723
box -33 -37 33 37
use M2M3_PR  M2M3_PR_61
timestamp 1626908933
transform 1 0 13680 0 1 7723
box -33 -37 33 37
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_68
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_187
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_68
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_187
timestamp 1626908933
transform 1 0 13700 0 1 7992
box -100 -49 100 49
use L1M1_PR  L1M1_PR_944
timestamp 1626908933
transform 1 0 13584 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_547
timestamp 1626908933
transform 1 0 13488 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_442
timestamp 1626908933
transform 1 0 13584 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_45
timestamp 1626908933
transform 1 0 13488 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_196
timestamp 1626908933
transform 1 0 13728 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_83
timestamp 1626908933
transform 1 0 13728 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_116
timestamp 1626908933
transform 1 0 13632 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_34
timestamp 1626908933
transform 1 0 13632 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_132
timestamp 1626908933
transform 1 0 13920 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_302
timestamp 1626908933
transform 1 0 13920 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_40
timestamp 1626908933
transform 1 0 0 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_210
timestamp 1626908933
transform 1 0 0 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_386
timestamp 1626908933
transform 1 0 240 0 1 8843
box -32 -32 32 32
use M1M2_PR  M1M2_PR_851
timestamp 1626908933
transform 1 0 240 0 1 8843
box -32 -32 32 32
use M2M3_PR  M2M3_PR_34
timestamp 1626908933
transform 1 0 240 0 1 8943
box -33 -37 33 37
use M2M3_PR  M2M3_PR_76
timestamp 1626908933
transform 1 0 240 0 1 8943
box -33 -37 33 37
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_59
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_178
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_59
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_178
timestamp 1626908933
transform 1 0 500 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_96
timestamp 1626908933
transform 1 0 96 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_199
timestamp 1626908933
transform 1 0 96 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_209
timestamp 1626908933
transform 1 0 1248 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_39
timestamp 1626908933
transform 1 0 1248 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_227
timestamp 1626908933
transform 1 0 864 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_107
timestamp 1626908933
transform 1 0 864 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_183
timestamp 1626908933
transform 1 0 1344 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_80
timestamp 1626908933
transform 1 0 1344 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_33
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_115
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_90
timestamp 1626908933
transform 1 0 2112 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_210
timestamp 1626908933
transform 1 0 2112 0 -1 9324
box -38 -49 422 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_167
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_48
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_167
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_48
timestamp 1626908933
transform 1 0 2900 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_524
timestamp 1626908933
transform 1 0 2736 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_22
timestamp 1626908933
transform 1 0 2736 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_671
timestamp 1626908933
transform 1 0 2832 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_206
timestamp 1626908933
transform 1 0 2832 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_762
timestamp 1626908933
transform 1 0 2928 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_260
timestamp 1626908933
transform 1 0 2928 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_24
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_56
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 710 715
use L1M1_PR  L1M1_PR_993
timestamp 1626908933
transform 1 0 3024 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_841
timestamp 1626908933
transform 1 0 3024 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_491
timestamp 1626908933
transform 1 0 3024 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_339
timestamp 1626908933
transform 1 0 3024 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_914
timestamp 1626908933
transform 1 0 3024 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_912
timestamp 1626908933
transform 1 0 3120 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_449
timestamp 1626908933
transform 1 0 3024 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_447
timestamp 1626908933
transform 1 0 3120 0 1 8399
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_208
timestamp 1626908933
transform 1 0 3264 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_38
timestamp 1626908933
transform 1 0 3264 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_202
timestamp 1626908933
transform 1 0 3360 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_82
timestamp 1626908933
transform 1 0 3360 0 -1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_282
timestamp 1626908933
transform 1 0 3888 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_283
timestamp 1626908933
transform 1 0 3888 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_322
timestamp 1626908933
transform 1 0 3600 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_747
timestamp 1626908933
transform 1 0 3888 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_748
timestamp 1626908933
transform 1 0 3888 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_787
timestamp 1626908933
transform 1 0 3600 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_378
timestamp 1626908933
transform 1 0 3792 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_880
timestamp 1626908933
transform 1 0 3792 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_64
timestamp 1626908933
transform 1 0 3744 0 -1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_27
timestamp 1626908933
transform 1 0 3744 0 -1 9324
box -38 -49 1958 715
use L1M1_PR  L1M1_PR_840
timestamp 1626908933
transform 1 0 4176 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_338
timestamp 1626908933
transform 1 0 4176 0 1 8991
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_156
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_37
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_156
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_37
timestamp 1626908933
transform 1 0 5300 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_523
timestamp 1626908933
transform 1 0 5328 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_21
timestamp 1626908933
transform 1 0 5328 0 1 8917
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_185
timestamp 1626908933
transform 1 0 5664 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_65
timestamp 1626908933
transform 1 0 5664 0 -1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_620
timestamp 1626908933
transform 1 0 6288 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_118
timestamp 1626908933
transform 1 0 6288 0 1 8399
box -29 -23 29 23
use M1M2_PR  M1M2_PR_582
timestamp 1626908933
transform 1 0 6192 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_117
timestamp 1626908933
transform 1 0 6192 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_522
timestamp 1626908933
transform 1 0 6096 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_20
timestamp 1626908933
transform 1 0 6096 0 1 8917
box -29 -23 29 23
use M1M2_PR  M1M2_PR_810
timestamp 1626908933
transform 1 0 6288 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_345
timestamp 1626908933
transform 1 0 6288 0 1 9065
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_197
timestamp 1626908933
transform 1 0 6048 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_84
timestamp 1626908933
transform 1 0 6048 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_46
timestamp 1626908933
transform 1 0 6240 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_17
timestamp 1626908933
transform 1 0 6240 0 -1 9324
box -38 -49 326 715
use L1M1_PR  L1M1_PR_903
timestamp 1626908933
transform 1 0 6480 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_692
timestamp 1626908933
transform 1 0 6384 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_401
timestamp 1626908933
transform 1 0 6480 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_190
timestamp 1626908933
transform 1 0 6384 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_623
timestamp 1626908933
transform 1 0 6672 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_158
timestamp 1626908933
transform 1 0 6672 0 1 8769
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_303
timestamp 1626908933
transform 1 0 6720 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_133
timestamp 1626908933
transform 1 0 6720 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_198
timestamp 1626908933
transform 1 0 6528 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_85
timestamp 1626908933
transform 1 0 6528 0 -1 9324
box -38 -49 230 715
use L1M1_PR  L1M1_PR_181
timestamp 1626908933
transform 1 0 7056 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_683
timestamp 1626908933
transform 1 0 7056 0 1 8769
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_32
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_114
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_66
timestamp 1626908933
transform 1 0 7344 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_531
timestamp 1626908933
transform 1 0 7344 0 1 8769
box -32 -32 32 32
use L1M1_PR  L1M1_PR_189
timestamp 1626908933
transform 1 0 7152 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_192
timestamp 1626908933
transform 1 0 7248 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_691
timestamp 1626908933
transform 1 0 7152 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_694
timestamp 1626908933
transform 1 0 7248 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_20
timestamp 1626908933
transform -1 0 7488 0 -1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_54
timestamp 1626908933
transform -1 0 7488 0 -1 9324
box -38 -49 710 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_145
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_26
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_145
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_26
timestamp 1626908933
transform 1 0 7700 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_568
timestamp 1626908933
transform 1 0 7728 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_66
timestamp 1626908933
transform 1 0 7728 0 1 8769
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_199
timestamp 1626908933
transform 1 0 7584 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_86
timestamp 1626908933
transform 1 0 7584 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_45
timestamp 1626908933
transform 1 0 7776 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_16
timestamp 1626908933
transform 1 0 7776 0 -1 9324
box -38 -49 326 715
use L1M1_PR  L1M1_PR_141
timestamp 1626908933
transform 1 0 7920 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_191
timestamp 1626908933
transform 1 0 7920 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_643
timestamp 1626908933
transform 1 0 7920 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_693
timestamp 1626908933
transform 1 0 7920 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_87
timestamp 1626908933
transform 1 0 8064 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_200
timestamp 1626908933
transform 1 0 8064 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_134
timestamp 1626908933
transform 1 0 8256 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_304
timestamp 1626908933
transform 1 0 8256 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_135
timestamp 1626908933
transform 1 0 8112 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_600
timestamp 1626908933
transform 1 0 8112 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_416
timestamp 1626908933
transform 1 0 8112 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_918
timestamp 1626908933
transform 1 0 8112 0 1 9139
box -29 -23 29 23
use L1M1_PR  L1M1_PR_652
timestamp 1626908933
transform 1 0 8688 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_150
timestamp 1626908933
transform 1 0 8688 0 1 8399
box -29 -23 29 23
use M1M2_PR  M1M2_PR_604
timestamp 1626908933
transform 1 0 8784 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_139
timestamp 1626908933
transform 1 0 8784 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_656
timestamp 1626908933
transform 1 0 8688 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_651
timestamp 1626908933
transform 1 0 8784 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_154
timestamp 1626908933
transform 1 0 8688 0 1 8917
box -29 -23 29 23
use L1M1_PR  L1M1_PR_149
timestamp 1626908933
transform 1 0 8784 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_603
timestamp 1626908933
transform 1 0 8784 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_138
timestamp 1626908933
transform 1 0 8784 0 1 8769
box -32 -32 32 32
use L1M1_PR  L1M1_PR_653
timestamp 1626908933
transform 1 0 8688 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_151
timestamp 1626908933
transform 1 0 8688 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_10
timestamp 1626908933
transform 1 0 8352 0 -1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_44
timestamp 1626908933
transform 1 0 8352 0 -1 9324
box -38 -49 710 715
use M1M2_PR  M1M2_PR_608
timestamp 1626908933
transform 1 0 9360 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_605
timestamp 1626908933
transform 1 0 9072 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_517
timestamp 1626908933
transform 1 0 9936 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_143
timestamp 1626908933
transform 1 0 9360 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_140
timestamp 1626908933
transform 1 0 9072 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_52
timestamp 1626908933
transform 1 0 9936 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_131
timestamp 1626908933
transform 1 0 9024 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_28
timestamp 1626908933
transform 1 0 9024 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_40
timestamp 1626908933
transform -1 0 11712 0 -1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_3
timestamp 1626908933
transform -1 0 11712 0 -1 9324
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_134
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_15
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_134
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_15
timestamp 1626908933
transform 1 0 10100 0 1 8658
box -100 -49 100 49
use L1M1_PR  L1M1_PR_917
timestamp 1626908933
transform 1 0 10416 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_415
timestamp 1626908933
transform 1 0 10416 0 1 8399
box -29 -23 29 23
use M1M2_PR  M1M2_PR_828
timestamp 1626908933
transform 1 0 10704 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_363
timestamp 1626908933
transform 1 0 10704 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_50
timestamp 1626908933
transform 1 0 11088 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_552
timestamp 1626908933
transform 1 0 11088 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_267
timestamp 1626908933
transform 1 0 11472 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_732
timestamp 1626908933
transform 1 0 11472 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_191
timestamp 1626908933
transform 1 0 11088 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_656
timestamp 1626908933
transform 1 0 11088 0 1 8917
box -32 -32 32 32
use L1M1_PR  L1M1_PR_319
timestamp 1626908933
transform 1 0 11280 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_821
timestamp 1626908933
transform 1 0 11280 0 1 9065
box -29 -23 29 23
use M1M2_PR  M1M2_PR_298
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_763
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_355
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_857
timestamp 1626908933
transform 1 0 11664 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_118
timestamp 1626908933
transform 1 0 11712 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_15
timestamp 1626908933
transform 1 0 11712 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_31
timestamp 1626908933
transform 1 0 12480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_113
timestamp 1626908933
transform 1 0 12480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_135
timestamp 1626908933
transform 1 0 12576 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_305
timestamp 1626908933
transform 1 0 12576 0 -1 9324
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_4
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_123
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_4
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_123
timestamp 1626908933
transform 1 0 12500 0 1 8658
box -100 -49 100 49
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_15
timestamp 1626908933
transform 1 0 12672 0 -1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_47
timestamp 1626908933
transform 1 0 12672 0 -1 9324
box -38 -49 710 715
use M1M2_PR  M1M2_PR_49
timestamp 1626908933
transform 1 0 12912 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_423
timestamp 1626908933
transform 1 0 12912 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_424
timestamp 1626908933
transform 1 0 12912 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_514
timestamp 1626908933
transform 1 0 12912 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_888
timestamp 1626908933
transform 1 0 12912 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_889
timestamp 1626908933
transform 1 0 12912 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_49
timestamp 1626908933
transform 1 0 12816 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_551
timestamp 1626908933
transform 1 0 12816 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_238
timestamp 1626908933
transform 1 0 13008 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_320
timestamp 1626908933
transform 1 0 13008 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_463
timestamp 1626908933
transform 1 0 13104 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_740
timestamp 1626908933
transform 1 0 13008 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_822
timestamp 1626908933
transform 1 0 13008 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_965
timestamp 1626908933
transform 1 0 13104 0 1 8991
box -29 -23 29 23
use M2M3_PR  M2M3_PR_17
timestamp 1626908933
transform 1 0 13008 0 1 8943
box -33 -37 33 37
use M2M3_PR  M2M3_PR_59
timestamp 1626908933
transform 1 0 13008 0 1 8943
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_88
timestamp 1626908933
transform 1 0 13344 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_201
timestamp 1626908933
transform 1 0 13344 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_45
timestamp 1626908933
transform 1 0 13392 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_510
timestamp 1626908933
transform 1 0 13392 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_318
timestamp 1626908933
transform 1 0 13296 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_820
timestamp 1626908933
transform 1 0 13296 0 1 9065
box -29 -23 29 23
use M1M2_PR  M1M2_PR_651
timestamp 1626908933
transform 1 0 13488 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_186
timestamp 1626908933
transform 1 0 13488 0 1 8769
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_306
timestamp 1626908933
transform 1 0 13536 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_136
timestamp 1626908933
transform 1 0 13536 0 -1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_735
timestamp 1626908933
transform 1 0 13776 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_546
timestamp 1626908933
transform 1 0 13680 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_233
timestamp 1626908933
transform 1 0 13776 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_44
timestamp 1626908933
transform 1 0 13680 0 1 9065
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_57
timestamp 1626908933
transform 1 0 13632 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_28
timestamp 1626908933
transform 1 0 13632 0 -1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_137
timestamp 1626908933
transform 1 0 13920 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_307
timestamp 1626908933
transform 1 0 13920 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_353
timestamp 1626908933
transform 1 0 13968 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_818
timestamp 1626908933
transform 1 0 13968 0 1 9065
box -32 -32 32 32
use L1M1_PR  L1M1_PR_409
timestamp 1626908933
transform 1 0 13872 0 1 9065
box -29 -23 29 23
use L1M1_PR  L1M1_PR_911
timestamp 1626908933
transform 1 0 13872 0 1 9065
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_308
timestamp 1626908933
transform 1 0 192 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_138
timestamp 1626908933
transform 1 0 192 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_852
timestamp 1626908933
transform 1 0 240 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_387
timestamp 1626908933
transform 1 0 240 0 1 9435
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_207
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_37
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_112
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_30
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_202
timestamp 1626908933
transform 1 0 0 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_89
timestamp 1626908933
transform 1 0 0 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_86
timestamp 1626908933
transform 1 0 480 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_189
timestamp 1626908933
transform 1 0 480 0 1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_435
timestamp 1626908933
transform 1 0 1296 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_937
timestamp 1626908933
transform 1 0 1296 0 1 9435
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_112
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_231
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_112
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_231
timestamp 1626908933
transform 1 0 1700 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_214
timestamp 1626908933
transform 1 0 1680 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_679
timestamp 1626908933
transform 1 0 1680 0 1 9805
box -32 -32 32 32
use L1M1_PR  L1M1_PR_25
timestamp 1626908933
transform 1 0 1392 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_266
timestamp 1626908933
transform 1 0 1584 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_497
timestamp 1626908933
transform 1 0 1680 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_527
timestamp 1626908933
transform 1 0 1392 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_768
timestamp 1626908933
transform 1 0 1584 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_999
timestamp 1626908933
transform 1 0 1680 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_23
timestamp 1626908933
transform 1 0 1248 0 1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_55
timestamp 1626908933
transform 1 0 1248 0 1 9324
box -38 -49 710 715
use L1M1_PR  L1M1_PR_837
timestamp 1626908933
transform 1 0 1872 0 1 9805
box -29 -23 29 23
use L1M1_PR  L1M1_PR_335
timestamp 1626908933
transform 1 0 1872 0 1 9805
box -29 -23 29 23
use M1M2_PR  M1M2_PR_922
timestamp 1626908933
transform 1 0 1872 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_457
timestamp 1626908933
transform 1 0 1872 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_217
timestamp 1626908933
transform 1 0 1920 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_97
timestamp 1626908933
transform 1 0 1920 0 1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_9
timestamp 1626908933
transform 1 0 2352 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_474
timestamp 1626908933
transform 1 0 2352 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_8
timestamp 1626908933
transform 1 0 2352 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_510
timestamp 1626908933
transform 1 0 2352 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_279
timestamp 1626908933
transform 1 0 2352 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_744
timestamp 1626908933
transform 1 0 2352 0 1 9805
box -32 -32 32 32
use L1M1_PR  L1M1_PR_122
timestamp 1626908933
transform 1 0 2448 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_624
timestamp 1626908933
transform 1 0 2448 0 1 9731
box -29 -23 29 23
use M1M2_PR  M1M2_PR_341
timestamp 1626908933
transform 1 0 2160 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_806
timestamp 1626908933
transform 1 0 2160 0 1 9879
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_29
timestamp 1626908933
transform 1 0 2304 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_0
timestamp 1626908933
transform 1 0 2304 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_86
timestamp 1626908933
transform 1 0 2688 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_206
timestamp 1626908933
transform 1 0 2688 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_36
timestamp 1626908933
transform 1 0 2592 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_206
timestamp 1626908933
transform 1 0 2592 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_397
timestamp 1626908933
transform 1 0 2640 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_434
timestamp 1626908933
transform 1 0 2640 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_899
timestamp 1626908933
transform 1 0 2640 0 1 9879
box -29 -23 29 23
use L1M1_PR  L1M1_PR_936
timestamp 1626908933
transform 1 0 2640 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_281
timestamp 1626908933
transform 1 0 3408 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_746
timestamp 1626908933
transform 1 0 3408 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_337
timestamp 1626908933
transform 1 0 3216 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_839
timestamp 1626908933
transform 1 0 3216 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_448
timestamp 1626908933
transform 1 0 3024 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_913
timestamp 1626908933
transform 1 0 3024 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_280
timestamp 1626908933
transform 1 0 3408 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_745
timestamp 1626908933
transform 1 0 3408 0 1 9509
box -32 -32 32 32
use L1M1_PR  L1M1_PR_336
timestamp 1626908933
transform 1 0 3504 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_838
timestamp 1626908933
transform 1 0 3504 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_382
timestamp 1626908933
transform 1 0 3120 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_884
timestamp 1626908933
transform 1 0 3120 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_321
timestamp 1626908933
transform 1 0 3600 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_786
timestamp 1626908933
transform 1 0 3600 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_147
timestamp 1626908933
transform 1 0 3120 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_612
timestamp 1626908933
transform 1 0 3120 0 1 9879
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_63
timestamp 1626908933
transform 1 0 3072 0 1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_26
timestamp 1626908933
transform 1 0 3072 0 1 9324
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_221
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_102
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_221
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_102
timestamp 1626908933
transform 1 0 4100 0 1 9324
box -100 -49 100 49
use L1M1_PR  L1M1_PR_526
timestamp 1626908933
transform 1 0 4656 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_24
timestamp 1626908933
transform 1 0 4656 0 1 9435
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_205
timestamp 1626908933
transform 1 0 5280 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_35
timestamp 1626908933
transform 1 0 5280 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_130
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_17
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_152
timestamp 1626908933
transform 1 0 5376 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_49
timestamp 1626908933
transform 1 0 5376 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_111
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_29
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_116
timestamp 1626908933
transform 1 0 6192 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_581
timestamp 1626908933
transform 1 0 6192 0 1 9435
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_92
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_211
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_92
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_211
timestamp 1626908933
transform 1 0 6500 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_119
timestamp 1626908933
transform 1 0 6576 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_584
timestamp 1626908933
transform 1 0 6576 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_120
timestamp 1626908933
transform 1 0 6480 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_121
timestamp 1626908933
transform 1 0 6480 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_622
timestamp 1626908933
transform 1 0 6480 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_623
timestamp 1626908933
transform 1 0 6480 0 1 9731
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_2
timestamp 1626908933
transform 1 0 6144 0 1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_36
timestamp 1626908933
transform 1 0 6144 0 1 9324
box -38 -49 710 715
use L1M1_PR  L1M1_PR_619
timestamp 1626908933
transform 1 0 6768 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_117
timestamp 1626908933
transform 1 0 6768 0 1 9435
box -29 -23 29 23
use M1M2_PR  M1M2_PR_831
timestamp 1626908933
transform 1 0 6960 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_366
timestamp 1626908933
transform 1 0 6960 0 1 9509
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_309
timestamp 1626908933
transform 1 0 7008 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_139
timestamp 1626908933
transform 1 0 7008 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_203
timestamp 1626908933
transform 1 0 6816 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_90
timestamp 1626908933
transform 1 0 6816 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_34
timestamp 1626908933
transform 1 0 7104 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_5
timestamp 1626908933
transform 1 0 7104 0 1 9324
box -38 -49 326 715
use L1M1_PR  L1M1_PR_904
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_646
timestamp 1626908933
transform 1 0 7248 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_525
timestamp 1626908933
transform 1 0 7152 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_402
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_144
timestamp 1626908933
transform 1 0 7248 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_23
timestamp 1626908933
transform 1 0 7152 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_811
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_346
timestamp 1626908933
transform 1 0 7344 0 1 9583
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_204
timestamp 1626908933
transform 1 0 7392 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_91
timestamp 1626908933
transform 1 0 7392 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_42
timestamp 1626908933
transform -1 0 8352 0 1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_8
timestamp 1626908933
transform -1 0 8352 0 1 9324
box -38 -49 710 715
use L1M1_PR  L1M1_PR_644
timestamp 1626908933
transform 1 0 7728 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_142
timestamp 1626908933
transform 1 0 7728 0 1 9435
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_310
timestamp 1626908933
transform 1 0 7584 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_140
timestamp 1626908933
transform 1 0 7584 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_16
timestamp 1626908933
transform 1 0 8352 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_129
timestamp 1626908933
transform 1 0 8352 0 1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_134
timestamp 1626908933
transform 1 0 8112 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_599
timestamp 1626908933
transform 1 0 8112 0 1 9435
box -32 -32 32 32
use L1M1_PR  L1M1_PR_143
timestamp 1626908933
transform 1 0 8016 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_146
timestamp 1626908933
transform 1 0 8016 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_645
timestamp 1626908933
transform 1 0 8016 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_648
timestamp 1626908933
transform 1 0 8016 0 1 9731
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_48
timestamp 1626908933
transform 1 0 8544 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_168
timestamp 1626908933
transform 1 0 8544 0 1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_142
timestamp 1626908933
transform 1 0 9360 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_607
timestamp 1626908933
transform 1 0 9360 0 1 9435
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_82
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_201
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_82
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_201
timestamp 1626908933
transform 1 0 8900 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_144
timestamp 1626908933
transform 1 0 8976 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_145
timestamp 1626908933
transform 1 0 8976 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_609
timestamp 1626908933
transform 1 0 8976 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_610
timestamp 1626908933
transform 1 0 8976 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_156
timestamp 1626908933
transform 1 0 9264 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_157
timestamp 1626908933
transform 1 0 9168 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_658
timestamp 1626908933
transform 1 0 9264 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_659
timestamp 1626908933
transform 1 0 9168 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_11
timestamp 1626908933
transform 1 0 8928 0 1 9324
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_45
timestamp 1626908933
transform 1 0 8928 0 1 9324
box -38 -49 710 715
use L1M1_PR  L1M1_PR_655
timestamp 1626908933
transform 1 0 9552 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_153
timestamp 1626908933
transform 1 0 9552 0 1 9435
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_161
timestamp 1626908933
transform 1 0 9600 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_41
timestamp 1626908933
transform 1 0 9600 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_110
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_28
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_554
timestamp 1626908933
transform 1 0 10128 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_52
timestamp 1626908933
transform 1 0 10128 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_516
timestamp 1626908933
transform 1 0 10128 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_515
timestamp 1626908933
transform 1 0 10128 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_51
timestamp 1626908933
transform 1 0 10128 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_50
timestamp 1626908933
transform 1 0 10128 0 1 9583
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_311
timestamp 1626908933
transform 1 0 10080 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_141
timestamp 1626908933
transform 1 0 10080 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_657
timestamp 1626908933
transform 1 0 10320 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_553
timestamp 1626908933
transform 1 0 10224 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_155
timestamp 1626908933
transform 1 0 10320 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_51
timestamp 1626908933
transform 1 0 10224 0 1 9583
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_36
timestamp 1626908933
transform 1 0 10176 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_7
timestamp 1626908933
transform 1 0 10176 0 1 9324
box -38 -49 326 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_4
timestamp 1626908933
transform 1 0 10464 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_11
timestamp 1626908933
transform 1 0 10464 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_92
timestamp 1626908933
transform 1 0 10848 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_205
timestamp 1626908933
transform 1 0 10848 0 1 9324
box -38 -49 230 715
use L1M1_PR  L1M1_PR_411
timestamp 1626908933
transform 1 0 10512 0 1 9731
box -29 -23 29 23
use L1M1_PR  L1M1_PR_913
timestamp 1626908933
transform 1 0 10512 0 1 9731
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_142
timestamp 1626908933
transform 1 0 11040 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_312
timestamp 1626908933
transform 1 0 11040 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_358
timestamp 1626908933
transform 1 0 11184 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_860
timestamp 1626908933
transform 1 0 11184 0 1 9657
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_72
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_191
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_72
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_191
timestamp 1626908933
transform 1 0 11300 0 1 9324
box -100 -49 100 49
use M1M2_PR  M1M2_PR_266
timestamp 1626908933
transform 1 0 11472 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_731
timestamp 1626908933
transform 1 0 11472 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_321
timestamp 1626908933
transform 1 0 11568 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_823
timestamp 1626908933
transform 1 0 11568 0 1 9583
box -29 -23 29 23
use M1M2_PR  M1M2_PR_297
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_762
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_55
timestamp 1626908933
transform 1 0 11136 0 1 9324
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_18
timestamp 1626908933
transform 1 0 11136 0 1 9324
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_401
timestamp 1626908933
transform 1 0 12720 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_866
timestamp 1626908933
transform 1 0 12720 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_443
timestamp 1626908933
transform 1 0 12720 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_945
timestamp 1626908933
transform 1 0 12720 0 1 9213
box -29 -23 29 23
use M1M2_PR  M1M2_PR_365
timestamp 1626908933
transform 1 0 12720 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_830
timestamp 1626908933
transform 1 0 12720 0 1 9509
box -32 -32 32 32
use M2M3_PR  M2M3_PR_16
timestamp 1626908933
transform 1 0 12720 0 1 9553
box -33 -37 33 37
use M2M3_PR  M2M3_PR_58
timestamp 1626908933
transform 1 0 12720 0 1 9553
box -33 -37 33 37
use M1M2_PR  M1M2_PR_355
timestamp 1626908933
transform 1 0 12816 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_820
timestamp 1626908933
transform 1 0 12816 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_137
timestamp 1626908933
transform 1 0 12720 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_602
timestamp 1626908933
transform 1 0 12720 0 1 9879
box -32 -32 32 32
use L1M1_PR  L1M1_PR_550
timestamp 1626908933
transform 1 0 12912 0 1 9435
box -29 -23 29 23
use L1M1_PR  L1M1_PR_48
timestamp 1626908933
transform 1 0 12912 0 1 9435
box -29 -23 29 23
use M1M2_PR  M1M2_PR_513
timestamp 1626908933
transform 1 0 12912 0 1 9435
box -32 -32 32 32
use M1M2_PR  M1M2_PR_48
timestamp 1626908933
transform 1 0 12912 0 1 9435
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_124
timestamp 1626908933
transform 1 0 13056 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_4
timestamp 1626908933
transform 1 0 13056 0 1 9324
box -38 -49 422 715
use M1M2_PR  M1M2_PR_364
timestamp 1626908933
transform 1 0 13488 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_829
timestamp 1626908933
transform 1 0 13488 0 1 9213
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_27
timestamp 1626908933
transform 1 0 13632 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_109
timestamp 1626908933
transform 1 0 13632 0 1 9324
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_67
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_186
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_67
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_186
timestamp 1626908933
transform 1 0 13700 0 1 9324
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_93
timestamp 1626908933
transform 1 0 13440 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_94
timestamp 1626908933
transform 1 0 13728 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_206
timestamp 1626908933
transform 1 0 13440 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_207
timestamp 1626908933
transform 1 0 13728 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_313
timestamp 1626908933
transform 1 0 13920 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_143
timestamp 1626908933
transform 1 0 13920 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_318
timestamp 1626908933
transform 1 0 192 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_204
timestamp 1626908933
transform 1 0 0 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_148
timestamp 1626908933
transform 1 0 192 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_34
timestamp 1626908933
transform 1 0 0 0 -1 10656
box -38 -49 134 715
use M2M3_PR  M2M3_PR_77
timestamp 1626908933
transform 1 0 240 0 1 10041
box -33 -37 33 37
use M2M3_PR  M2M3_PR_35
timestamp 1626908933
transform 1 0 240 0 1 10041
box -33 -37 33 37
use M1M2_PR  M1M2_PR_853
timestamp 1626908933
transform 1 0 240 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_388
timestamp 1626908933
transform 1 0 240 0 1 10545
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_105
timestamp 1626908933
transform 1 0 288 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_23
timestamp 1626908933
transform 1 0 288 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_210
timestamp 1626908933
transform 1 0 0 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_97
timestamp 1626908933
transform 1 0 0 0 1 10656
box -38 -49 230 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_58
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_177
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_58
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_177
timestamp 1626908933
transform 1 0 500 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_85
timestamp 1626908933
transform 1 0 768 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_95
timestamp 1626908933
transform 1 0 96 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_188
timestamp 1626908933
transform 1 0 768 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_198
timestamp 1626908933
transform 1 0 96 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_114
timestamp 1626908933
transform 1 0 384 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_234
timestamp 1626908933
transform 1 0 384 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_15
timestamp 1626908933
transform 1 0 864 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_128
timestamp 1626908933
transform 1 0 864 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_33
timestamp 1626908933
transform 1 0 1056 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_203
timestamp 1626908933
transform 1 0 1056 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_436
timestamp 1626908933
transform 1 0 1200 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_938
timestamp 1626908933
transform 1 0 1200 0 1 10545
box -29 -23 29 23
use M1M2_PR  M1M2_PR_678
timestamp 1626908933
transform 1 0 1680 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_213
timestamp 1626908933
transform 1 0 1680 0 1 10175
box -32 -32 32 32
use L1M1_PR  L1M1_PR_530
timestamp 1626908933
transform 1 0 1296 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_28
timestamp 1626908933
transform 1 0 1296 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_491
timestamp 1626908933
transform 1 0 1296 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_26
timestamp 1626908933
transform 1 0 1296 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1000
timestamp 1626908933
transform 1 0 1584 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_769
timestamp 1626908933
transform 1 0 1488 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_498
timestamp 1626908933
transform 1 0 1584 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_267
timestamp 1626908933
transform 1 0 1488 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_478
timestamp 1626908933
transform 1 0 1680 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_13
timestamp 1626908933
transform 1 0 1680 0 1 10397
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_230
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_111
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_230
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_111
timestamp 1626908933
transform 1 0 1700 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_74
timestamp 1626908933
transform 1 0 1536 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_177
timestamp 1626908933
transform 1 0 1536 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_22
timestamp 1626908933
transform 1 0 1152 0 -1 10656
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_54
timestamp 1626908933
transform 1 0 1152 0 -1 10656
box -38 -49 710 715
use L1M1_PR  L1M1_PR_835
timestamp 1626908933
transform 1 0 1776 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_333
timestamp 1626908933
transform 1 0 1776 0 1 10545
box -29 -23 29 23
use M1M2_PR  M1M2_PR_921
timestamp 1626908933
transform 1 0 1872 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_456
timestamp 1626908933
transform 1 0 1872 0 1 10249
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_202
timestamp 1626908933
transform 1 0 1824 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_32
timestamp 1626908933
transform 1 0 1824 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_216
timestamp 1626908933
transform 1 0 1920 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_96
timestamp 1626908933
transform 1 0 1920 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_31
timestamp 1626908933
transform 1 0 2304 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_201
timestamp 1626908933
transform 1 0 2304 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_26
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_108
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_95
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_208
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_144
timestamp 1626908933
transform 1 0 2400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_314
timestamp 1626908933
transform 1 0 2400 0 -1 10656
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_166
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_47
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_166
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_47
timestamp 1626908933
transform 1 0 2900 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_660
timestamp 1626908933
transform 1 0 2928 0 1 10175
box -29 -23 29 23
use L1M1_PR  L1M1_PR_158
timestamp 1626908933
transform 1 0 2928 0 1 10175
box -29 -23 29 23
use M1M2_PR  M1M2_PR_916
timestamp 1626908933
transform 1 0 2832 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_451
timestamp 1626908933
transform 1 0 2832 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_514
timestamp 1626908933
transform 1 0 2832 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_12
timestamp 1626908933
transform 1 0 2832 0 1 10397
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_35
timestamp 1626908933
transform 1 0 2784 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_6
timestamp 1626908933
transform 1 0 2784 0 -1 10656
box -38 -49 326 715
use L1M1_PR  L1M1_PR_900
timestamp 1626908933
transform 1 0 3120 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_398
timestamp 1626908933
transform 1 0 3120 0 1 10545
box -29 -23 29 23
use M1M2_PR  M1M2_PR_807
timestamp 1626908933
transform 1 0 3216 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_611
timestamp 1626908933
transform 1 0 3120 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_342
timestamp 1626908933
transform 1 0 3216 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_146
timestamp 1626908933
transform 1 0 3120 0 1 10175
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_315
timestamp 1626908933
transform 1 0 3456 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_145
timestamp 1626908933
transform 1 0 3456 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_12
timestamp 1626908933
transform 1 0 3072 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_5
timestamp 1626908933
transform 1 0 3072 0 -1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_320
timestamp 1626908933
transform 1 0 3600 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_785
timestamp 1626908933
transform 1 0 3600 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_380
timestamp 1626908933
transform 1 0 3600 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_882
timestamp 1626908933
transform 1 0 3600 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_332
timestamp 1626908933
transform 1 0 3984 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_834
timestamp 1626908933
transform 1 0 3984 0 1 10397
box -29 -23 29 23
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_62
timestamp 1626908933
transform -1 0 4224 0 1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_61
timestamp 1626908933
transform 1 0 3552 0 -1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_25
timestamp 1626908933
transform -1 0 4224 0 1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_24
timestamp 1626908933
transform 1 0 3552 0 -1 10656
box -38 -49 1958 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_220
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_101
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_220
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_101
timestamp 1626908933
transform 1 0 4100 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_160
timestamp 1626908933
transform 1 0 4224 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_57
timestamp 1626908933
transform 1 0 4224 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_104
timestamp 1626908933
transform 1 0 4992 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_22
timestamp 1626908933
transform 1 0 4992 0 1 10656
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_155
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_36
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_155
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_36
timestamp 1626908933
transform 1 0 5300 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_532
timestamp 1626908933
transform 1 0 5328 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_30
timestamp 1626908933
transform 1 0 5328 0 1 10545
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_319
timestamp 1626908933
transform 1 0 5280 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_200
timestamp 1626908933
transform 1 0 5472 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_149
timestamp 1626908933
transform 1 0 5280 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_30
timestamp 1626908933
transform 1 0 5472 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_211
timestamp 1626908933
transform 1 0 5088 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_98
timestamp 1626908933
transform 1 0 5088 0 1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_27
timestamp 1626908933
transform 1 0 5520 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_492
timestamp 1626908933
transform 1 0 5520 0 1 10545
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_48
timestamp 1626908933
transform 1 0 5568 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_151
timestamp 1626908933
transform 1 0 5568 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_60
timestamp 1626908933
transform 1 0 5376 0 1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_23
timestamp 1626908933
transform 1 0 5376 0 1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_61
timestamp 1626908933
transform 1 0 6336 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_181
timestamp 1626908933
transform 1 0 6336 0 -1 10656
box -38 -49 422 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_91
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_210
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_91
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_210
timestamp 1626908933
transform 1 0 6500 0 1 10656
box -100 -49 100 49
use M1M2_PR  M1M2_PR_118
timestamp 1626908933
transform 1 0 6576 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_583
timestamp 1626908933
transform 1 0 6576 0 1 10101
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_41
timestamp 1626908933
transform 1 0 6720 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_144
timestamp 1626908933
transform 1 0 6720 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_25
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_107
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_99
timestamp 1626908933
transform 1 0 7296 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_212
timestamp 1626908933
transform 1 0 7296 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_150
timestamp 1626908933
transform 1 0 7488 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_320
timestamp 1626908933
transform 1 0 7488 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_315
timestamp 1626908933
transform 1 0 7632 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_780
timestamp 1626908933
transform 1 0 7632 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_368
timestamp 1626908933
transform 1 0 7632 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_870
timestamp 1626908933
transform 1 0 7632 0 1 10323
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_25
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_144
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_25
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_144
timestamp 1626908933
transform 1 0 7700 0 1 9990
box -100 -49 100 49
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_59
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_58
timestamp 1626908933
transform 1 0 7584 0 1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_22
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_21
timestamp 1626908933
transform 1 0 7584 0 1 10656
box -38 -49 1958 715
use M1M2_PR  M1M2_PR_275
timestamp 1626908933
transform 1 0 8016 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_740
timestamp 1626908933
transform 1 0 8016 0 1 10397
box -32 -32 32 32
use L1M1_PR  L1M1_PR_328
timestamp 1626908933
transform 1 0 8016 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_830
timestamp 1626908933
transform 1 0 8016 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_36
timestamp 1626908933
transform 1 0 8592 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_501
timestamp 1626908933
transform 1 0 8592 0 1 10545
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_81
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_200
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_81
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_200
timestamp 1626908933
transform 1 0 8900 0 1 10656
box -100 -49 100 49
use L1M1_PR  L1M1_PR_35
timestamp 1626908933
transform 1 0 9168 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_537
timestamp 1626908933
transform 1 0 9168 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_865
timestamp 1626908933
transform 1 0 9648 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_363
timestamp 1626908933
transform 1 0 9648 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_736
timestamp 1626908933
transform 1 0 9456 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_271
timestamp 1626908933
transform 1 0 9456 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_316
timestamp 1626908933
transform 1 0 9504 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_199
timestamp 1626908933
transform 1 0 9504 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_146
timestamp 1626908933
transform 1 0 9504 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_29
timestamp 1626908933
transform 1 0 9504 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_160
timestamp 1626908933
transform 1 0 9600 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_40
timestamp 1626908933
transform 1 0 9600 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_21
timestamp 1626908933
transform 1 0 9984 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_103
timestamp 1626908933
transform 1 0 9984 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_57
timestamp 1626908933
transform 1 0 9600 0 -1 10656
box -38 -49 1958 715
use sky130_fd_sc_hs__dfxtp_4  sky130_fd_sc_hs__dfxtp_4_20
timestamp 1626908933
transform 1 0 9600 0 -1 10656
box -38 -49 1958 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_14
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_133
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_14
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_133
timestamp 1626908933
transform 1 0 10100 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_324
timestamp 1626908933
transform 1 0 10032 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_826
timestamp 1626908933
transform 1 0 10032 0 1 10397
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_23
timestamp 1626908933
transform 1 0 10464 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_126
timestamp 1626908933
transform 1 0 10464 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_34
timestamp 1626908933
transform 1 0 10080 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_154
timestamp 1626908933
transform 1 0 10080 0 1 10656
box -38 -49 422 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_71
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_190
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_71
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_190
timestamp 1626908933
transform 1 0 11300 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_28
timestamp 1626908933
transform 1 0 11616 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_198
timestamp 1626908933
transform 1 0 11616 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_43
timestamp 1626908933
transform 1 0 11376 0 1 10471
box -29 -23 29 23
use L1M1_PR  L1M1_PR_545
timestamp 1626908933
transform 1 0 11376 0 1 10471
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_18
timestamp 1626908933
transform 1 0 11520 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_24
timestamp 1626908933
transform 1 0 11232 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_138
timestamp 1626908933
transform 1 0 11520 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_144
timestamp 1626908933
transform 1 0 11232 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_209
timestamp 1626908933
transform 1 0 11904 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_96
timestamp 1626908933
transform 1 0 11904 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_117
timestamp 1626908933
transform 1 0 11712 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_14
timestamp 1626908933
transform 1 0 11712 0 1 10656
box -38 -49 806 715
use L1M1_PR  L1M1_PR_544
timestamp 1626908933
transform 1 0 12144 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_42
timestamp 1626908933
transform 1 0 12144 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_621
timestamp 1626908933
transform 1 0 12240 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_119
timestamp 1626908933
transform 1 0 12240 0 1 10101
box -29 -23 29 23
use M1M2_PR  M1M2_PR_508
timestamp 1626908933
transform 1 0 12336 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_43
timestamp 1626908933
transform 1 0 12336 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_317
timestamp 1626908933
transform 1 0 12384 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_147
timestamp 1626908933
transform 1 0 12384 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_30
timestamp 1626908933
transform 1 0 12096 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_1
timestamp 1626908933
transform 1 0 12096 0 -1 10656
box -38 -49 326 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_122
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_3
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_122
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_3
timestamp 1626908933
transform 1 0 12500 0 1 9990
box -100 -49 100 49
use L1M1_PR  L1M1_PR_910
timestamp 1626908933
transform 1 0 12432 0 1 10545
box -29 -23 29 23
use L1M1_PR  L1M1_PR_408
timestamp 1626908933
transform 1 0 12432 0 1 10545
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_106
timestamp 1626908933
transform 1 0 12480 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_24
timestamp 1626908933
transform 1 0 12480 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_601
timestamp 1626908933
transform 1 0 12720 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_136
timestamp 1626908933
transform 1 0 12720 0 1 10101
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_10
timestamp 1626908933
transform 1 0 12480 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_11
timestamp 1626908933
transform 1 0 12576 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_130
timestamp 1626908933
transform 1 0 12480 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_131
timestamp 1626908933
transform 1 0 12576 0 -1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_647
timestamp 1626908933
transform 1 0 13104 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_145
timestamp 1626908933
transform 1 0 13104 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_912
timestamp 1626908933
transform 1 0 13200 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_549
timestamp 1626908933
transform 1 0 13008 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_410
timestamp 1626908933
transform 1 0 13200 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_47
timestamp 1626908933
transform 1 0 13008 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_512
timestamp 1626908933
transform 1 0 12912 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_47
timestamp 1626908933
transform 1 0 12912 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_127
timestamp 1626908933
transform 1 0 13248 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_14
timestamp 1626908933
transform 1 0 13248 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_33
timestamp 1626908933
transform 1 0 12960 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_4
timestamp 1626908933
transform 1 0 12960 0 -1 10656
box -38 -49 326 715
use M1M2_PR  M1M2_PR_819
timestamp 1626908933
transform 1 0 13296 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_354
timestamp 1626908933
transform 1 0 13296 0 1 10397
box -32 -32 32 32
use M2M3_PR  M2M3_PR_15
timestamp 1626908933
transform 1 0 13584 0 1 10285
box -33 -37 33 37
use M2M3_PR  M2M3_PR_57
timestamp 1626908933
transform 1 0 13584 0 1 10285
box -33 -37 33 37
use M1M2_PR  M1M2_PR_352
timestamp 1626908933
transform 1 0 13488 0 1 10545
box -32 -32 32 32
use M1M2_PR  M1M2_PR_817
timestamp 1626908933
transform 1 0 13488 0 1 10545
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_66
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_185
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_66
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_185
timestamp 1626908933
transform 1 0 13700 0 1 10656
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_20
timestamp 1626908933
transform 1 0 13632 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_102
timestamp 1626908933
transform 1 0 13632 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_4
timestamp 1626908933
transform 1 0 12864 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_107
timestamp 1626908933
transform 1 0 12864 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1
timestamp 1626908933
transform 1 0 13440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_121
timestamp 1626908933
transform 1 0 13440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_321
timestamp 1626908933
transform 1 0 13920 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_151
timestamp 1626908933
transform 1 0 13920 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_213
timestamp 1626908933
transform 1 0 13728 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_126
timestamp 1626908933
transform 1 0 13824 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_100
timestamp 1626908933
transform 1 0 13728 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_13
timestamp 1626908933
transform 1 0 13824 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_27
timestamp 1626908933
transform 1 0 0 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_197
timestamp 1626908933
transform 1 0 0 0 -1 11988
box -38 -49 134 715
use M2M3_PR  M2M3_PR_36
timestamp 1626908933
transform 1 0 240 0 1 11139
box -33 -37 33 37
use M2M3_PR  M2M3_PR_78
timestamp 1626908933
transform 1 0 240 0 1 11139
box -33 -37 33 37
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_57
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_176
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_57
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_176
timestamp 1626908933
transform 1 0 500 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_94
timestamp 1626908933
transform 1 0 96 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_197
timestamp 1626908933
transform 1 0 96 0 -1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_490
timestamp 1626908933
transform 1 0 1296 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_25
timestamp 1626908933
transform 1 0 1296 0 1 10767
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_196
timestamp 1626908933
transform 1 0 1248 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_26
timestamp 1626908933
transform 1 0 1248 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_226
timestamp 1626908933
transform 1 0 864 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_106
timestamp 1626908933
transform 1 0 864 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_182
timestamp 1626908933
transform 1 0 1344 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_79
timestamp 1626908933
transform 1 0 1344 0 -1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_278
timestamp 1626908933
transform 1 0 2352 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_743
timestamp 1626908933
transform 1 0 2352 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_529
timestamp 1626908933
transform 1 0 2448 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_27
timestamp 1626908933
transform 1 0 2448 0 1 10767
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_101
timestamp 1626908933
transform 1 0 2496 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_19
timestamp 1626908933
transform 1 0 2496 0 -1 11988
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_165
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_46
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_165
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_46
timestamp 1626908933
transform 1 0 2900 0 1 11322
box -100 -49 100 49
use M1M2_PR  M1M2_PR_915
timestamp 1626908933
transform 1 0 2832 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_450
timestamp 1626908933
transform 1 0 2832 0 1 11211
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_68
timestamp 1626908933
transform 1 0 2592 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_171
timestamp 1626908933
transform 1 0 2592 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_89
timestamp 1626908933
transform 1 0 2112 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_209
timestamp 1626908933
transform 1 0 2112 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_784
timestamp 1626908933
transform 1 0 3600 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_319
timestamp 1626908933
transform 1 0 3600 0 1 10989
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_201
timestamp 1626908933
transform 1 0 3360 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_81
timestamp 1626908933
transform 1 0 3360 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_836
timestamp 1626908933
transform 1 0 3792 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_334
timestamp 1626908933
transform 1 0 3792 0 1 10915
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_163
timestamp 1626908933
transform 1 0 3744 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_60
timestamp 1626908933
transform 1 0 3744 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_53
timestamp 1626908933
transform 1 0 4608 0 -1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_21
timestamp 1626908933
transform 1 0 4608 0 -1 11988
box -38 -49 710 715
use L1M1_PR  L1M1_PR_879
timestamp 1626908933
transform 1 0 4176 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_377
timestamp 1626908933
transform 1 0 4176 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_322
timestamp 1626908933
transform 1 0 4512 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_152
timestamp 1626908933
transform 1 0 4512 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_489
timestamp 1626908933
transform 1 0 4848 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_24
timestamp 1626908933
transform 1 0 4848 0 1 10767
box -32 -32 32 32
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_154
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_35
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_154
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_35
timestamp 1626908933
transform 1 0 5300 0 1 11322
box -100 -49 100 49
use M1M2_PR  M1M2_PR_909
timestamp 1626908933
transform 1 0 5136 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_444
timestamp 1626908933
transform 1 0 5136 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_833
timestamp 1626908933
transform 1 0 5232 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_331
timestamp 1626908933
transform 1 0 5232 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_12
timestamp 1626908933
transform 1 0 5280 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_125
timestamp 1626908933
transform 1 0 5280 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_25
timestamp 1626908933
transform 1 0 5472 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_195
timestamp 1626908933
transform 1 0 5472 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_374
timestamp 1626908933
transform 1 0 5424 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_876
timestamp 1626908933
transform 1 0 5424 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_47
timestamp 1626908933
transform 1 0 5568 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_150
timestamp 1626908933
transform 1 0 5568 0 -1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_832
timestamp 1626908933
transform 1 0 5808 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_330
timestamp 1626908933
transform 1 0 5808 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_742
timestamp 1626908933
transform 1 0 5808 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_741
timestamp 1626908933
transform 1 0 5808 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_277
timestamp 1626908933
transform 1 0 5808 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_276
timestamp 1626908933
transform 1 0 5808 0 1 11433
box -32 -32 32 32
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_52
timestamp 1626908933
transform 1 0 6336 0 -1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_20
timestamp 1626908933
transform 1 0 6336 0 -1 11988
box -38 -49 710 715
use M1M2_PR  M1M2_PR_498
timestamp 1626908933
transform 1 0 6576 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_33
timestamp 1626908933
transform 1 0 6576 0 1 11211
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_24
timestamp 1626908933
transform 1 0 7008 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_194
timestamp 1626908933
transform 1 0 7008 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_33
timestamp 1626908933
transform 1 0 6960 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_329
timestamp 1626908933
transform 1 0 6960 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_535
timestamp 1626908933
transform 1 0 6960 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_831
timestamp 1626908933
transform 1 0 6960 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_18
timestamp 1626908933
transform 1 0 7488 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_100
timestamp 1626908933
transform 1 0 7488 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_56
timestamp 1626908933
transform 1 0 7104 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_176
timestamp 1626908933
transform 1 0 7104 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_314
timestamp 1626908933
transform 1 0 7632 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_779
timestamp 1626908933
transform 1 0 7632 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_367
timestamp 1626908933
transform 1 0 7632 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_869
timestamp 1626908933
transform 1 0 7632 0 1 10989
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_24
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_143
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_24
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_143
timestamp 1626908933
transform 1 0 7700 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_19
timestamp 1626908933
transform 1 0 7584 0 -1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_51
timestamp 1626908933
transform 1 0 7584 0 -1 11988
box -38 -49 710 715
use M1M2_PR  M1M2_PR_273
timestamp 1626908933
transform 1 0 8208 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_738
timestamp 1626908933
transform 1 0 8208 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_327
timestamp 1626908933
transform 1 0 8016 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_829
timestamp 1626908933
transform 1 0 8016 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_272
timestamp 1626908933
transform 1 0 8208 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_274
timestamp 1626908933
transform 1 0 8016 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_737
timestamp 1626908933
transform 1 0 8208 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_739
timestamp 1626908933
transform 1 0 8016 0 1 11433
box -32 -32 32 32
use L1M1_PR  L1M1_PR_326
timestamp 1626908933
transform 1 0 8208 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_828
timestamp 1626908933
transform 1 0 8208 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_6
timestamp 1626908933
transform 1 0 8256 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_13
timestamp 1626908933
transform 1 0 8256 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_18
timestamp 1626908933
transform 1 0 8640 0 -1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__a22o_1  sky130_fd_sc_hs__a22o_1_50
timestamp 1626908933
transform 1 0 8640 0 -1 11988
box -38 -49 710 715
use M1M2_PR  M1M2_PR_506
timestamp 1626908933
transform 1 0 8784 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_41
timestamp 1626908933
transform 1 0 8784 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_540
timestamp 1626908933
transform 1 0 9168 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_38
timestamp 1626908933
transform 1 0 9168 0 1 11211
box -29 -23 29 23
use M1M2_PR  M1M2_PR_496
timestamp 1626908933
transform 1 0 9264 0 1 11137
box -32 -32 32 32
use M1M2_PR  M1M2_PR_31
timestamp 1626908933
transform 1 0 9264 0 1 11137
box -32 -32 32 32
use L1M1_PR  L1M1_PR_827
timestamp 1626908933
transform 1 0 9264 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_325
timestamp 1626908933
transform 1 0 9264 0 1 11433
box -29 -23 29 23
use M1M2_PR  M1M2_PR_735
timestamp 1626908933
transform 1 0 9456 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_270
timestamp 1626908933
transform 1 0 9456 0 1 11433
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_44
timestamp 1626908933
transform 1 0 9312 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_164
timestamp 1626908933
transform 1 0 9312 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_733
timestamp 1626908933
transform 1 0 9840 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_231
timestamp 1626908933
transform 1 0 9840 0 1 11433
box -29 -23 29 23
use M1M2_PR  M1M2_PR_649
timestamp 1626908933
transform 1 0 9648 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_184
timestamp 1626908933
transform 1 0 9648 0 1 11433
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_193
timestamp 1626908933
transform 1 0 9984 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_23
timestamp 1626908933
transform 1 0 9984 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_54
timestamp 1626908933
transform 1 0 9696 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_25
timestamp 1626908933
transform 1 0 9696 0 -1 11988
box -38 -49 326 715
use M1M2_PR  M1M2_PR_362
timestamp 1626908933
transform 1 0 10704 0 1 10841
box -32 -32 32 32
use M1M2_PR  M1M2_PR_827
timestamp 1626908933
transform 1 0 10704 0 1 10841
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_13
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_132
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_13
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_132
timestamp 1626908933
transform 1 0 10100 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_22
timestamp 1626908933
transform 1 0 10464 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_125
timestamp 1626908933
transform 1 0 10464 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_33
timestamp 1626908933
transform 1 0 10080 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_153
timestamp 1626908933
transform 1 0 10080 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_192
timestamp 1626908933
transform 1 0 11616 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_22
timestamp 1626908933
transform 1 0 11616 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_143
timestamp 1626908933
transform 1 0 11232 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_23
timestamp 1626908933
transform 1 0 11232 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_116
timestamp 1626908933
transform 1 0 11712 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_13
timestamp 1626908933
transform 1 0 11712 0 -1 11988
box -38 -49 806 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_121
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_2
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_121
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_2
timestamp 1626908933
transform 1 0 12500 0 1 11322
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_99
timestamp 1626908933
transform 1 0 12480 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_17
timestamp 1626908933
transform 1 0 12480 0 -1 11988
box -38 -49 134 715
use M2M3_PR  M2M3_PR_56
timestamp 1626908933
transform 1 0 12720 0 1 10895
box -33 -37 33 37
use M2M3_PR  M2M3_PR_14
timestamp 1626908933
transform 1 0 12720 0 1 10895
box -33 -37 33 37
use M1M2_PR  M1M2_PR_826
timestamp 1626908933
transform 1 0 12720 0 1 10841
box -32 -32 32 32
use M1M2_PR  M1M2_PR_361
timestamp 1626908933
transform 1 0 12720 0 1 10841
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_9
timestamp 1626908933
transform 1 0 12576 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_129
timestamp 1626908933
transform 1 0 12576 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_106
timestamp 1626908933
transform 1 0 12960 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_3
timestamp 1626908933
transform 1 0 12960 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_323
timestamp 1626908933
transform 1 0 13920 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_153
timestamp 1626908933
transform 1 0 13920 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_214
timestamp 1626908933
transform 1 0 13728 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_101
timestamp 1626908933
transform 1 0 13728 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_324
timestamp 1626908933
transform 1 0 192 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_154
timestamp 1626908933
transform 1 0 192 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_855
timestamp 1626908933
transform 1 0 240 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_854
timestamp 1626908933
transform 1 0 240 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_390
timestamp 1626908933
transform 1 0 240 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_389
timestamp 1626908933
transform 1 0 240 0 1 11729
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_98
timestamp 1626908933
transform 1 0 288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_16
timestamp 1626908933
transform 1 0 288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_215
timestamp 1626908933
transform 1 0 0 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_102
timestamp 1626908933
transform 1 0 0 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_84
timestamp 1626908933
transform 1 0 768 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_187
timestamp 1626908933
transform 1 0 768 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_113
timestamp 1626908933
transform 1 0 384 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_233
timestamp 1626908933
transform 1 0 384 0 1 11988
box -38 -49 422 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_229
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_110
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_229
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_110
timestamp 1626908933
transform 1 0 1700 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_220
timestamp 1626908933
transform 1 0 1536 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_100
timestamp 1626908933
transform 1 0 1536 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_675
timestamp 1626908933
transform 1 0 1872 0 1 11507
box -32 -32 32 32
use M1M2_PR  M1M2_PR_210
timestamp 1626908933
transform 1 0 1872 0 1 11507
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_176
timestamp 1626908933
transform 1 0 1920 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_73
timestamp 1626908933
transform 1 0 1920 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_20
timestamp 1626908933
transform 1 0 3552 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_49
timestamp 1626908933
transform 1 0 3552 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_64
timestamp 1626908933
transform 1 0 2784 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_167
timestamp 1626908933
transform 1 0 2784 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_103
timestamp 1626908933
transform 1 0 3840 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_216
timestamp 1626908933
transform 1 0 3840 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_21
timestamp 1626908933
transform 1 0 2688 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_191
timestamp 1626908933
transform 1 0 2688 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_155
timestamp 1626908933
transform 1 0 4032 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_325
timestamp 1626908933
transform 1 0 4032 0 1 11988
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_100
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_219
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_100
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_219
timestamp 1626908933
transform 1 0 4100 0 1 11988
box -100 -49 100 49
use L1M1_PR  L1M1_PR_31
timestamp 1626908933
transform 1 0 4560 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_437
timestamp 1626908933
transform 1 0 4464 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_533
timestamp 1626908933
transform 1 0 4560 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_939
timestamp 1626908933
transform 1 0 4464 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_24
timestamp 1626908933
transform 1 0 4128 0 1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_58
timestamp 1626908933
transform 1 0 4128 0 1 11988
box -38 -49 710 715
use L1M1_PR  L1M1_PR_987
timestamp 1626908933
transform 1 0 5040 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_756
timestamp 1626908933
transform 1 0 4944 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_485
timestamp 1626908933
transform 1 0 5040 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_254
timestamp 1626908933
transform 1 0 4944 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_97
timestamp 1626908933
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_15
timestamp 1626908933
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_218
timestamp 1626908933
transform 1 0 5088 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_217
timestamp 1626908933
transform 1 0 4800 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_105
timestamp 1626908933
transform 1 0 5088 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_104
timestamp 1626908933
transform 1 0 4800 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_21
timestamp 1626908933
transform 1 0 5376 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_50
timestamp 1626908933
transform 1 0 5376 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_156
timestamp 1626908933
transform 1 0 5280 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_326
timestamp 1626908933
transform 1 0 5280 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_29
timestamp 1626908933
transform 1 0 5424 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_443
timestamp 1626908933
transform 1 0 5232 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_494
timestamp 1626908933
transform 1 0 5424 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_908
timestamp 1626908933
transform 1 0 5232 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_57
timestamp 1626908933
transform 1 0 5952 0 1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_23
timestamp 1626908933
transform 1 0 5952 0 1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_327
timestamp 1626908933
transform 1 0 5856 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_157
timestamp 1626908933
transform 1 0 5856 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_219
timestamp 1626908933
transform 1 0 5664 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_106
timestamp 1626908933
transform 1 0 5664 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_438
timestamp 1626908933
transform 1 0 6384 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_940
timestamp 1626908933
transform 1 0 6384 0 1 11877
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_209
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_90
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_209
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_90
timestamp 1626908933
transform 1 0 6500 0 1 11988
box -100 -49 100 49
use L1M1_PR  L1M1_PR_536
timestamp 1626908933
transform 1 0 6480 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_34
timestamp 1626908933
transform 1 0 6480 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_497
timestamp 1626908933
transform 1 0 6576 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_32
timestamp 1626908933
transform 1 0 6576 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_984
timestamp 1626908933
transform 1 0 6768 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_754
timestamp 1626908933
transform 1 0 6672 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_482
timestamp 1626908933
transform 1 0 6768 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_252
timestamp 1626908933
transform 1 0 6672 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_328
timestamp 1626908933
transform 1 0 6624 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_158
timestamp 1626908933
transform 1 0 6624 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_22
timestamp 1626908933
transform 1 0 6720 0 1 11988
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_56
timestamp 1626908933
transform 1 0 6720 0 1 11988
box -38 -49 710 715
use M1M2_PR  M1M2_PR_120
timestamp 1626908933
transform 1 0 7056 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_392
timestamp 1626908933
transform 1 0 6864 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_585
timestamp 1626908933
transform 1 0 7056 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_857
timestamp 1626908933
transform 1 0 6864 0 1 11877
box -32 -32 32 32
use L1M1_PR  L1M1_PR_123
timestamp 1626908933
transform 1 0 7344 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_439
timestamp 1626908933
transform 1 0 7632 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_625
timestamp 1626908933
transform 1 0 7344 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_941
timestamp 1626908933
transform 1 0 7632 0 1 11877
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_37
timestamp 1626908933
transform 1 0 7392 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_140
timestamp 1626908933
transform 1 0 7392 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_749
timestamp 1626908933
transform 1 0 7920 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_539
timestamp 1626908933
transform 1 0 7728 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_247
timestamp 1626908933
transform 1 0 7920 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_37
timestamp 1626908933
transform 1 0 7728 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_503
timestamp 1626908933
transform 1 0 7728 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_502
timestamp 1626908933
transform 1 0 7728 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_38
timestamp 1626908933
transform 1 0 7728 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_37
timestamp 1626908933
transform 1 0 7728 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_20
timestamp 1626908933
transform 1 0 8160 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_190
timestamp 1626908933
transform 1 0 8160 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_395
timestamp 1626908933
transform 1 0 8400 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_860
timestamp 1626908933
transform 1 0 8400 0 1 11877
box -32 -32 32 32
use L1M1_PR  L1M1_PR_478
timestamp 1626908933
transform 1 0 8016 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_980
timestamp 1626908933
transform 1 0 8016 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_35
timestamp 1626908933
transform 1 0 8592 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_40
timestamp 1626908933
transform 1 0 8784 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_500
timestamp 1626908933
transform 1 0 8592 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_505
timestamp 1626908933
transform 1 0 8784 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_40
timestamp 1626908933
transform 1 0 8784 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_440
timestamp 1626908933
transform 1 0 8592 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_542
timestamp 1626908933
transform 1 0 8784 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_942
timestamp 1626908933
transform 1 0 8592 0 1 11877
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_31
timestamp 1626908933
transform 1 0 8640 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_134
timestamp 1626908933
transform 1 0 8640 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_50
timestamp 1626908933
transform 1 0 8256 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_170
timestamp 1626908933
transform 1 0 8256 0 1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_245
timestamp 1626908933
transform 1 0 8976 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_474
timestamp 1626908933
transform 1 0 9072 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_747
timestamp 1626908933
transform 1 0 8976 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_976
timestamp 1626908933
transform 1 0 9072 0 1 11655
box -29 -23 29 23
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_80
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_199
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_80
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_199
timestamp 1626908933
transform 1 0 8900 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_11
timestamp 1626908933
transform 1 0 9408 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_124
timestamp 1626908933
transform 1 0 9408 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_30
timestamp 1626908933
transform 1 0 9264 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_495
timestamp 1626908933
transform 1 0 9264 0 1 11729
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_39
timestamp 1626908933
transform 1 0 9600 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_159
timestamp 1626908933
transform 1 0 9600 0 1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_534
timestamp 1626908933
transform 1 0 9744 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_32
timestamp 1626908933
transform 1 0 9744 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_96
timestamp 1626908933
transform 1 0 9984 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_14
timestamp 1626908933
transform 1 0 9984 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_907
timestamp 1626908933
transform 1 0 10032 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_405
timestamp 1626908933
transform 1 0 10032 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_814
timestamp 1626908933
transform 1 0 10704 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_349
timestamp 1626908933
transform 1 0 10704 0 1 11877
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_152
timestamp 1626908933
transform 1 0 10080 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_32
timestamp 1626908933
transform 1 0 10080 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_124
timestamp 1626908933
transform 1 0 10464 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_21
timestamp 1626908933
transform 1 0 10464 0 1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_190
timestamp 1626908933
transform 1 0 11088 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_655
timestamp 1626908933
transform 1 0 11088 0 1 11581
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_70
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_189
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_70
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_189
timestamp 1626908933
transform 1 0 11300 0 1 11988
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_19
timestamp 1626908933
transform 1 0 11616 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_189
timestamp 1626908933
transform 1 0 11616 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_22
timestamp 1626908933
transform 1 0 11232 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_142
timestamp 1626908933
transform 1 0 11232 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_115
timestamp 1626908933
transform 1 0 11712 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_12
timestamp 1626908933
transform 1 0 11712 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_128
timestamp 1626908933
transform 1 0 12480 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_8
timestamp 1626908933
transform 1 0 12480 0 1 11988
box -38 -49 422 715
use M2M3_PR  M2M3_PR_13
timestamp 1626908933
transform 1 0 13008 0 1 11505
box -33 -37 33 37
use M2M3_PR  M2M3_PR_55
timestamp 1626908933
transform 1 0 13008 0 1 11505
box -33 -37 33 37
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_13
timestamp 1626908933
transform 1 0 13632 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_95
timestamp 1626908933
transform 1 0 13632 0 1 11988
box -38 -49 134 715
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_4
timestamp 1626908933
transform 1 0 13700 0 1 11965
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_12
timestamp 1626908933
transform 1 0 13700 0 1 11965
box -100 -26 100 26
use prbs_generator_syn_VIA11  prbs_generator_syn_VIA11_0
timestamp 1626908933
transform 1 0 13700 0 1 11952
box -100 -33 100 33
use prbs_generator_syn_VIA11  prbs_generator_syn_VIA11_1
timestamp 1626908933
transform 1 0 13700 0 1 11952
box -100 -33 100 33
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_2
timestamp 1626908933
transform 1 0 12864 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_105
timestamp 1626908933
transform 1 0 12864 0 1 11988
box -38 -49 806 715
use M2M3_PR  M2M3_PR_54
timestamp 1626908933
transform 1 0 13776 0 1 12115
box -33 -37 33 37
use M2M3_PR  M2M3_PR_12
timestamp 1626908933
transform 1 0 13776 0 1 12115
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_329
timestamp 1626908933
transform 1 0 13920 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_159
timestamp 1626908933
transform 1 0 13920 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_220
timestamp 1626908933
transform 1 0 13728 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_107
timestamp 1626908933
transform 1 0 13728 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_18
timestamp 1626908933
transform 1 0 0 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_188
timestamp 1626908933
transform 1 0 0 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_393
timestamp 1626908933
transform 1 0 240 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_858
timestamp 1626908933
transform 1 0 240 0 1 12987
box -32 -32 32 32
use M2M3_PR  M2M3_PR_37
timestamp 1626908933
transform 1 0 240 0 1 12237
box -33 -37 33 37
use M2M3_PR  M2M3_PR_79
timestamp 1626908933
transform 1 0 240 0 1 12237
box -33 -37 33 37
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_56
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_175
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_56
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_175
timestamp 1626908933
transform 1 0 500 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_93
timestamp 1626908933
transform 1 0 96 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_196
timestamp 1626908933
transform 1 0 96 0 -1 13320
box -38 -49 806 715
use M1M2_PR  M1M2_PR_481
timestamp 1626908933
transform 1 0 912 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_16
timestamp 1626908933
transform 1 0 912 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_187
timestamp 1626908933
transform 1 0 1248 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_17
timestamp 1626908933
transform 1 0 1248 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_225
timestamp 1626908933
transform 1 0 864 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_105
timestamp 1626908933
transform 1 0 864 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_181
timestamp 1626908933
transform 1 0 1344 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_78
timestamp 1626908933
transform 1 0 1344 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_12
timestamp 1626908933
transform 1 0 2496 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_94
timestamp 1626908933
transform 1 0 2496 0 -1 13320
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_45
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_164
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_45
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_164
timestamp 1626908933
transform 1 0 2900 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_67
timestamp 1626908933
transform 1 0 2592 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_170
timestamp 1626908933
transform 1 0 2592 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_88
timestamp 1626908933
transform 1 0 2112 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_208
timestamp 1626908933
transform 1 0 2112 0 -1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_516
timestamp 1626908933
transform 1 0 3504 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_14
timestamp 1626908933
transform 1 0 3504 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_200
timestamp 1626908933
transform 1 0 3360 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_80
timestamp 1626908933
transform 1 0 3360 0 -1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_901
timestamp 1626908933
transform 1 0 3792 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_710
timestamp 1626908933
transform 1 0 3696 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_399
timestamp 1626908933
transform 1 0 3792 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_208
timestamp 1626908933
transform 1 0 3696 0 1 12395
box -29 -23 29 23
use M1M2_PR  M1M2_PR_808
timestamp 1626908933
transform 1 0 3888 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_343
timestamp 1626908933
transform 1 0 3888 0 1 12247
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_162
timestamp 1626908933
transform 1 0 3744 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_59
timestamp 1626908933
transform 1 0 3744 0 -1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_709
timestamp 1626908933
transform 1 0 4464 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_708
timestamp 1626908933
transform 1 0 4464 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_207
timestamp 1626908933
transform 1 0 4464 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_206
timestamp 1626908933
transform 1 0 4464 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_191
timestamp 1626908933
transform 1 0 4512 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_71
timestamp 1626908933
transform 1 0 4512 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_330
timestamp 1626908933
transform 1 0 4896 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_160
timestamp 1626908933
transform 1 0 4896 0 -1 13320
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_153
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_34
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_153
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_34
timestamp 1626908933
transform 1 0 5300 0 1 12654
box -100 -49 100 49
use L1M1_PR  L1M1_PR_706
timestamp 1626908933
transform 1 0 5136 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_204
timestamp 1626908933
transform 1 0 5136 0 1 12395
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_51
timestamp 1626908933
transform 1 0 4992 0 -1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_22
timestamp 1626908933
transform 1 0 4992 0 -1 13320
box -38 -49 326 715
use L1M1_PR  L1M1_PR_531
timestamp 1626908933
transform 1 0 5424 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_29
timestamp 1626908933
transform 1 0 5424 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_493
timestamp 1626908933
transform 1 0 5424 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_28
timestamp 1626908933
transform 1 0 5424 0 1 12247
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_186
timestamp 1626908933
transform 1 0 5472 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_16
timestamp 1626908933
transform 1 0 5472 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_707
timestamp 1626908933
transform 1 0 5520 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_205
timestamp 1626908933
transform 1 0 5520 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_123
timestamp 1626908933
transform 1 0 5280 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_10
timestamp 1626908933
transform 1 0 5280 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_46
timestamp 1626908933
transform 1 0 5568 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_149
timestamp 1626908933
transform 1 0 5568 0 -1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_906
timestamp 1626908933
transform 1 0 5712 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_404
timestamp 1626908933
transform 1 0 5712 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_169
timestamp 1626908933
transform 1 0 6096 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_634
timestamp 1626908933
transform 1 0 6096 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_200
timestamp 1626908933
transform 1 0 6672 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_202
timestamp 1626908933
transform 1 0 6288 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_203
timestamp 1626908933
transform 1 0 6288 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_702
timestamp 1626908933
transform 1 0 6672 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_704
timestamp 1626908933
transform 1 0 6288 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_705
timestamp 1626908933
transform 1 0 6288 0 1 12395
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_40
timestamp 1626908933
transform 1 0 6720 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_143
timestamp 1626908933
transform 1 0 6720 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_60
timestamp 1626908933
transform 1 0 6336 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_180
timestamp 1626908933
transform 1 0 6336 0 -1 13320
box -38 -49 422 715
use M1M2_PR  M1M2_PR_391
timestamp 1626908933
transform 1 0 6864 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_856
timestamp 1626908933
transform 1 0 6864 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_198
timestamp 1626908933
transform 1 0 7056 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_199
timestamp 1626908933
transform 1 0 6960 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_700
timestamp 1626908933
transform 1 0 7056 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_701
timestamp 1626908933
transform 1 0 6960 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_167
timestamp 1626908933
transform 1 0 7536 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_632
timestamp 1626908933
transform 1 0 7536 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_166
timestamp 1626908933
transform 1 0 7536 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_631
timestamp 1626908933
transform 1 0 7536 0 1 12765
box -32 -32 32 32
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_23
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_142
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_23
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_142
timestamp 1626908933
transform 1 0 7700 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_11
timestamp 1626908933
transform 1 0 7488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_93
timestamp 1626908933
transform 1 0 7488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_26
timestamp 1626908933
transform -1 0 8256 0 -1 13320
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_60
timestamp 1626908933
transform -1 0 8256 0 -1 13320
box -38 -49 710 715
use L1M1_PR  L1M1_PR_718
timestamp 1626908933
transform 1 0 7920 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_699
timestamp 1626908933
transform 1 0 7824 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_216
timestamp 1626908933
transform 1 0 7920 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_197
timestamp 1626908933
transform 1 0 7824 0 1 12765
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_161
timestamp 1626908933
transform 1 0 8256 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_331
timestamp 1626908933
transform 1 0 8256 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_108
timestamp 1626908933
transform 1 0 8832 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_221
timestamp 1626908933
transform 1 0 8832 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_34
timestamp 1626908933
transform 1 0 8592 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_499
timestamp 1626908933
transform 1 0 8592 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_213
timestamp 1626908933
transform 1 0 8496 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_715
timestamp 1626908933
transform 1 0 8496 0 1 12913
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_3
timestamp 1626908933
transform 1 0 8352 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_0
timestamp 1626908933
transform 1 0 8352 0 -1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_717
timestamp 1626908933
transform 1 0 9168 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_215
timestamp 1626908933
transform 1 0 9168 0 1 12839
box -29 -23 29 23
use M1M2_PR  M1M2_PR_813
timestamp 1626908933
transform 1 0 9552 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_348
timestamp 1626908933
transform 1 0 9552 0 1 12543
box -32 -32 32 32
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_3
timestamp 1626908933
transform 1 0 9312 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_1
timestamp 1626908933
transform 1 0 9312 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_53
timestamp 1626908933
transform 1 0 9024 0 -1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_24
timestamp 1626908933
transform 1 0 9024 0 -1 13320
box -38 -49 326 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_131
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_12
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_131
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_12
timestamp 1626908933
transform 1 0 10100 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_151
timestamp 1626908933
transform 1 0 10080 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_31
timestamp 1626908933
transform 1 0 10080 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_123
timestamp 1626908933
transform 1 0 10464 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_20
timestamp 1626908933
transform 1 0 10464 0 -1 13320
box -38 -49 806 715
use M1M2_PR  M1M2_PR_822
timestamp 1626908933
transform 1 0 10896 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_357
timestamp 1626908933
transform 1 0 10896 0 1 12543
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_185
timestamp 1626908933
transform 1 0 11616 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_15
timestamp 1626908933
transform 1 0 11616 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_141
timestamp 1626908933
transform 1 0 11232 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_21
timestamp 1626908933
transform 1 0 11232 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_114
timestamp 1626908933
transform 1 0 11712 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_11
timestamp 1626908933
transform 1 0 11712 0 -1 13320
box -38 -49 806 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_120
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_1
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_120
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_1
timestamp 1626908933
transform 1 0 12500 0 1 12654
box -100 -49 100 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_92
timestamp 1626908933
transform 1 0 12480 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_10
timestamp 1626908933
transform 1 0 12480 0 -1 13320
box -38 -49 134 715
use M2M3_PR  M2M3_PR_53
timestamp 1626908933
transform 1 0 12720 0 1 12725
box -33 -37 33 37
use M2M3_PR  M2M3_PR_11
timestamp 1626908933
transform 1 0 12720 0 1 12725
box -33 -37 33 37
use M1M2_PR  M1M2_PR_821
timestamp 1626908933
transform 1 0 12720 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_816
timestamp 1626908933
transform 1 0 12720 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_356
timestamp 1626908933
transform 1 0 12720 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_351
timestamp 1626908933
transform 1 0 12720 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_7
timestamp 1626908933
transform 1 0 12576 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_127
timestamp 1626908933
transform 1 0 12576 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_104
timestamp 1626908933
transform 1 0 12960 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1
timestamp 1626908933
transform 1 0 12960 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_332
timestamp 1626908933
transform 1 0 13920 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_162
timestamp 1626908933
transform 1 0 13920 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_222
timestamp 1626908933
transform 1 0 13728 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_109
timestamp 1626908933
transform 1 0 13728 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_9
timestamp 1626908933
transform 1 0 288 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_91
timestamp 1626908933
transform 1 0 288 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_110
timestamp 1626908933
transform 1 0 0 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_223
timestamp 1626908933
transform 1 0 0 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_163
timestamp 1626908933
transform 1 0 192 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_333
timestamp 1626908933
transform 1 0 192 0 1 13320
box -38 -49 134 715
use M2M3_PR  M2M3_PR_38
timestamp 1626908933
transform 1 0 240 0 1 13335
box -33 -37 33 37
use M2M3_PR  M2M3_PR_80
timestamp 1626908933
transform 1 0 240 0 1 13335
box -33 -37 33 37
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_83
timestamp 1626908933
transform 1 0 768 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_186
timestamp 1626908933
transform 1 0 768 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_112
timestamp 1626908933
transform 1 0 384 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_232
timestamp 1626908933
transform 1 0 384 0 1 13320
box -38 -49 422 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_228
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_109
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_228
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_109
timestamp 1626908933
transform 1 0 1700 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_219
timestamp 1626908933
transform 1 0 1536 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_99
timestamp 1626908933
transform 1 0 1536 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_175
timestamp 1626908933
transform 1 0 1920 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_72
timestamp 1626908933
transform 1 0 1920 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_63
timestamp 1626908933
transform 1 0 3168 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_166
timestamp 1626908933
transform 1 0 3168 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_85
timestamp 1626908933
transform 1 0 2688 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_205
timestamp 1626908933
transform 1 0 2688 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_9
timestamp 1626908933
transform 1 0 3936 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_122
timestamp 1626908933
transform 1 0 3936 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_14
timestamp 1626908933
transform 1 0 3072 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_184
timestamp 1626908933
transform 1 0 3072 0 1 13320
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_218
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_99
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_218
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_99
timestamp 1626908933
transform 1 0 4100 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_183
timestamp 1626908933
transform 1 0 4128 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_13
timestamp 1626908933
transform 1 0 4128 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_159
timestamp 1626908933
transform 1 0 4224 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_56
timestamp 1626908933
transform 1 0 4224 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_90
timestamp 1626908933
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_8
timestamp 1626908933
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_520
timestamp 1626908933
transform 1 0 5040 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_18
timestamp 1626908933
transform 1 0 5040 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_484
timestamp 1626908933
transform 1 0 5040 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_19
timestamp 1626908933
transform 1 0 5040 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_902
timestamp 1626908933
transform 1 0 5232 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_714
timestamp 1626908933
transform 1 0 5232 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_400
timestamp 1626908933
transform 1 0 5232 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_212
timestamp 1626908933
transform 1 0 5232 0 1 13209
box -29 -23 29 23
use M1M2_PR  M1M2_PR_809
timestamp 1626908933
transform 1 0 5232 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_344
timestamp 1626908933
transform 1 0 5232 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_172
timestamp 1626908933
transform 1 0 5424 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_173
timestamp 1626908933
transform 1 0 5424 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_637
timestamp 1626908933
transform 1 0 5424 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_638
timestamp 1626908933
transform 1 0 5424 0 1 13209
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_45
timestamp 1626908933
transform 1 0 5088 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_148
timestamp 1626908933
transform 1 0 5088 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_59
timestamp 1626908933
transform 1 0 5856 0 1 13320
box -38 -49 710 715
use sky130_fd_sc_hs__xnor2_1  sky130_fd_sc_hs__xnor2_1_25
timestamp 1626908933
transform 1 0 5856 0 1 13320
box -38 -49 710 715
use M1M2_PR  M1M2_PR_168
timestamp 1626908933
transform 1 0 6096 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_171
timestamp 1626908933
transform 1 0 6096 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_633
timestamp 1626908933
transform 1 0 6096 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_636
timestamp 1626908933
transform 1 0 6096 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_209
timestamp 1626908933
transform 1 0 6192 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_211
timestamp 1626908933
transform 1 0 6192 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_711
timestamp 1626908933
transform 1 0 6192 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_713
timestamp 1626908933
transform 1 0 6192 0 1 13727
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_208
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_89
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_208
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_89
timestamp 1626908933
transform 1 0 6500 0 1 13320
box -100 -49 100 49
use L1M1_PR  L1M1_PR_703
timestamp 1626908933
transform 1 0 6480 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_201
timestamp 1626908933
transform 1 0 6480 0 1 13431
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_182
timestamp 1626908933
transform 1 0 6720 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_12
timestamp 1626908933
transform 1 0 6720 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_121
timestamp 1626908933
transform 1 0 6528 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_8
timestamp 1626908933
transform 1 0 6528 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_39
timestamp 1626908933
transform 1 0 6816 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_142
timestamp 1626908933
transform 1 0 6816 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_181
timestamp 1626908933
transform 1 0 7584 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_11
timestamp 1626908933
transform 1 0 7584 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_172
timestamp 1626908933
transform 1 0 7680 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_52
timestamp 1626908933
transform 1 0 7680 0 1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_716
timestamp 1626908933
transform 1 0 7920 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_214
timestamp 1626908933
transform 1 0 7920 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_908
timestamp 1626908933
transform 1 0 8688 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_538
timestamp 1626908933
transform 1 0 8592 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_406
timestamp 1626908933
transform 1 0 8688 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_36
timestamp 1626908933
transform 1 0 8592 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_165
timestamp 1626908933
transform 1 0 8832 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_45
timestamp 1626908933
transform 1 0 8832 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_136
timestamp 1626908933
transform 1 0 8064 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_33
timestamp 1626908933
transform 1 0 8064 0 1 13320
box -38 -49 806 715
use L1M1_PR  L1M1_PR_541
timestamp 1626908933
transform 1 0 9072 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_39
timestamp 1626908933
transform 1 0 9072 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_504
timestamp 1626908933
transform 1 0 9072 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_39
timestamp 1626908933
transform 1 0 9072 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_909
timestamp 1626908933
transform 1 0 9360 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_407
timestamp 1626908933
transform 1 0 9360 0 1 12987
box -29 -23 29 23
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_198
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_79
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_198
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_79
timestamp 1626908933
transform 1 0 8900 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_27
timestamp 1626908933
transform 1 0 9216 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_130
timestamp 1626908933
transform 1 0 9216 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_89
timestamp 1626908933
transform 1 0 9984 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_7
timestamp 1626908933
transform 1 0 9984 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_150
timestamp 1626908933
transform 1 0 10080 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_30
timestamp 1626908933
transform 1 0 10080 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_122
timestamp 1626908933
transform 1 0 10464 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_19
timestamp 1626908933
transform 1 0 10464 0 1 13320
box -38 -49 806 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_69
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_188
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_69
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_188
timestamp 1626908933
transform 1 0 11300 0 1 13320
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_10
timestamp 1626908933
transform 1 0 11616 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_180
timestamp 1626908933
transform 1 0 11616 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_350
timestamp 1626908933
transform 1 0 11664 0 1 13135
box -32 -32 32 32
use M1M2_PR  M1M2_PR_815
timestamp 1626908933
transform 1 0 11664 0 1 13135
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_20
timestamp 1626908933
transform 1 0 11232 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_140
timestamp 1626908933
transform 1 0 11232 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_113
timestamp 1626908933
transform 1 0 11712 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_10
timestamp 1626908933
transform 1 0 11712 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_126
timestamp 1626908933
transform 1 0 12480 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_6
timestamp 1626908933
transform 1 0 12480 0 1 13320
box -38 -49 422 715
use M2M3_PR  M2M3_PR_52
timestamp 1626908933
transform 1 0 13008 0 1 13335
box -33 -37 33 37
use M2M3_PR  M2M3_PR_10
timestamp 1626908933
transform 1 0 13008 0 1 13335
box -33 -37 33 37
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_103
timestamp 1626908933
transform 1 0 12864 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_0
timestamp 1626908933
transform 1 0 12864 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_88
timestamp 1626908933
transform 1 0 13632 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_6
timestamp 1626908933
transform 1 0 13632 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_334
timestamp 1626908933
transform 1 0 13920 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_164
timestamp 1626908933
transform 1 0 13920 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_224
timestamp 1626908933
transform 1 0 13728 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_111
timestamp 1626908933
transform 1 0 13728 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_165
timestamp 1626908933
transform 1 0 192 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_335
timestamp 1626908933
transform 1 0 192 0 -1 14652
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_174
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_55
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_174
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_55
timestamp 1626908933
transform 1 0 500 0 1 13986
box -100 -49 100 49
use M1M2_PR  M1M2_PR_861
timestamp 1626908933
transform 1 0 240 0 1 14171
box -32 -32 32 32
use M1M2_PR  M1M2_PR_396
timestamp 1626908933
transform 1 0 240 0 1 14171
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_179
timestamp 1626908933
transform 1 0 384 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_9
timestamp 1626908933
transform 1 0 384 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_87
timestamp 1626908933
transform 1 0 288 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_5
timestamp 1626908933
transform 1 0 288 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_112
timestamp 1626908933
transform 1 0 0 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_225
timestamp 1626908933
transform 1 0 0 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_231
timestamp 1626908933
transform 1 0 480 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_224
timestamp 1626908933
transform 1 0 864 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_111
timestamp 1626908933
transform 1 0 480 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_104
timestamp 1626908933
transform 1 0 864 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_223
timestamp 1626908933
transform 1 0 1248 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_103
timestamp 1626908933
transform 1 0 1248 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_218
timestamp 1626908933
transform 1 0 1632 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_98
timestamp 1626908933
transform 1 0 1632 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_178
timestamp 1626908933
transform 1 0 2016 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_8
timestamp 1626908933
transform 1 0 2016 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_207
timestamp 1626908933
transform 1 0 2112 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_87
timestamp 1626908933
transform 1 0 2112 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_4
timestamp 1626908933
transform 1 0 2496 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_86
timestamp 1626908933
transform 1 0 2496 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_7
timestamp 1626908933
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_177
timestamp 1626908933
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_44
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_163
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_44
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_163
timestamp 1626908933
transform 1 0 2900 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_84
timestamp 1626908933
transform 1 0 2688 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_204
timestamp 1626908933
transform 1 0 2688 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_203
timestamp 1626908933
transform 1 0 3072 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_83
timestamp 1626908933
transform 1 0 3072 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_199
timestamp 1626908933
transform 1 0 3456 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_195
timestamp 1626908933
transform 1 0 3840 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_79
timestamp 1626908933
transform 1 0 3456 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_75
timestamp 1626908933
transform 1 0 3840 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_194
timestamp 1626908933
transform 1 0 4224 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_74
timestamp 1626908933
transform 1 0 4224 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_488
timestamp 1626908933
transform 1 0 4848 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_23
timestamp 1626908933
transform 1 0 4848 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_189
timestamp 1626908933
transform 1 0 4608 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_69
timestamp 1626908933
transform 1 0 4608 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1626908933
transform 1 0 4992 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_85
timestamp 1626908933
transform 1 0 4992 0 -1 14652
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_33
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_152
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_33
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_152
timestamp 1626908933
transform 1 0 5300 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_67
timestamp 1626908933
transform 1 0 5280 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_187
timestamp 1626908933
transform 1 0 5280 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_7
timestamp 1626908933
transform 1 0 5088 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_120
timestamp 1626908933
transform 1 0 5088 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_119
timestamp 1626908933
transform 1 0 5664 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_6
timestamp 1626908933
transform 1 0 5664 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_336
timestamp 1626908933
transform 1 0 5856 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_166
timestamp 1626908933
transform 1 0 5856 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_52
timestamp 1626908933
transform 1 0 5952 0 -1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_23
timestamp 1626908933
transform 1 0 5952 0 -1 14652
box -38 -49 326 715
use M1M2_PR  M1M2_PR_170
timestamp 1626908933
transform 1 0 6096 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_635
timestamp 1626908933
transform 1 0 6096 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_210
timestamp 1626908933
transform 1 0 6096 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_712
timestamp 1626908933
transform 1 0 6096 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_26
timestamp 1626908933
transform 1 0 6000 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_403
timestamp 1626908933
transform 1 0 6192 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_528
timestamp 1626908933
transform 1 0 6000 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_905
timestamp 1626908933
transform 1 0 6192 0 1 14393
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_59
timestamp 1626908933
transform 1 0 6432 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_179
timestamp 1626908933
transform 1 0 6432 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_5
timestamp 1626908933
transform 1 0 6240 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_118
timestamp 1626908933
transform 1 0 6240 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_117
timestamp 1626908933
transform 1 0 6816 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_4
timestamp 1626908933
transform 1 0 6816 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_176
timestamp 1626908933
transform 1 0 7008 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_6
timestamp 1626908933
transform 1 0 7008 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_175
timestamp 1626908933
transform 1 0 7104 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_55
timestamp 1626908933
transform 1 0 7104 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1626908933
transform 1 0 7488 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_84
timestamp 1626908933
transform 1 0 7488 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_5
timestamp 1626908933
transform 1 0 7776 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_175
timestamp 1626908933
transform 1 0 7776 0 -1 14652
box -38 -49 134 715
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_22
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_141
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_22
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_141
timestamp 1626908933
transform 1 0 7700 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_3
timestamp 1626908933
transform 1 0 7584 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_116
timestamp 1626908933
transform 1 0 7584 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_171
timestamp 1626908933
transform 1 0 7872 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_51
timestamp 1626908933
transform 1 0 7872 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_859
timestamp 1626908933
transform 1 0 8400 0 1 14171
box -32 -32 32 32
use M1M2_PR  M1M2_PR_394
timestamp 1626908933
transform 1 0 8400 0 1 14171
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_169
timestamp 1626908933
transform 1 0 8256 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_49
timestamp 1626908933
transform 1 0 8256 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_812
timestamp 1626908933
transform 1 0 8592 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_347
timestamp 1626908933
transform 1 0 8592 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_167
timestamp 1626908933
transform 1 0 8640 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_47
timestamp 1626908933
transform 1 0 8640 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_174
timestamp 1626908933
transform 1 0 9216 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_4
timestamp 1626908933
transform 1 0 9216 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_115
timestamp 1626908933
transform 1 0 9024 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_2
timestamp 1626908933
transform 1 0 9024 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_163
timestamp 1626908933
transform 1 0 9312 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_43
timestamp 1626908933
transform 1 0 9312 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_114
timestamp 1626908933
transform 1 0 9696 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1
timestamp 1626908933
transform 1 0 9696 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_337
timestamp 1626908933
transform 1 0 9888 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_167
timestamp 1626908933
transform 1 0 9888 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_83
timestamp 1626908933
transform 1 0 9984 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1626908933
transform 1 0 9984 0 -1 14652
box -38 -49 134 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_130
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_11
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_130
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_11
timestamp 1626908933
transform 1 0 10100 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_149
timestamp 1626908933
transform 1 0 10080 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_29
timestamp 1626908933
transform 1 0 10080 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_148
timestamp 1626908933
transform 1 0 10464 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_146
timestamp 1626908933
transform 1 0 10848 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_28
timestamp 1626908933
transform 1 0 10464 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_26
timestamp 1626908933
transform 1 0 10848 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_139
timestamp 1626908933
transform 1 0 11232 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_19
timestamp 1626908933
transform 1 0 11232 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_173
timestamp 1626908933
transform 1 0 11808 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_3
timestamp 1626908933
transform 1 0 11808 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_113
timestamp 1626908933
transform 1 0 11616 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_0
timestamp 1626908933
transform 1 0 11616 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_136
timestamp 1626908933
transform 1 0 11904 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_16
timestamp 1626908933
transform 1 0 11904 0 -1 14652
box -38 -49 422 715
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_119
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA1  prbs_generator_syn_VIA1_0
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_119
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use prbs_generator_syn_VIA0  prbs_generator_syn_VIA0_0
timestamp 1626908933
transform 1 0 12500 0 1 13986
box -100 -49 100 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_338
timestamp 1626908933
transform 1 0 12384 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_172
timestamp 1626908933
transform 1 0 12288 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_168
timestamp 1626908933
transform 1 0 12384 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_2
timestamp 1626908933
transform 1 0 12288 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_171
timestamp 1626908933
transform 1 0 12576 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1
timestamp 1626908933
transform 1 0 12576 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_125
timestamp 1626908933
transform 1 0 12672 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_5
timestamp 1626908933
transform 1 0 12672 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_82
timestamp 1626908933
transform 1 0 12480 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0
timestamp 1626908933
transform 1 0 12480 0 -1 14652
box -38 -49 134 715
use M2M3_PR  M2M3_PR_51
timestamp 1626908933
transform 1 0 13200 0 1 13945
box -33 -37 33 37
use M2M3_PR  M2M3_PR_9
timestamp 1626908933
transform 1 0 13200 0 1 13945
box -33 -37 33 37
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_123
timestamp 1626908933
transform 1 0 13056 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_3
timestamp 1626908933
transform 1 0 13056 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_170
timestamp 1626908933
transform 1 0 13824 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_0
timestamp 1626908933
transform 1 0 13824 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_120
timestamp 1626908933
transform 1 0 13440 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_0
timestamp 1626908933
transform 1 0 13440 0 -1 14652
box -38 -49 422 715
use M2M3_PR  M2M3_PR_50
timestamp 1626908933
transform 1 0 13968 0 1 14189
box -33 -37 33 37
use M2M3_PR  M2M3_PR_8
timestamp 1626908933
transform 1 0 13968 0 1 14189
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_339
timestamp 1626908933
transform 1 0 13920 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_169
timestamp 1626908933
transform 1 0 13920 0 -1 14652
box -38 -49 134 715
use M2M3_PR  M2M3_PR_39
timestamp 1626908933
transform 1 0 240 0 1 14555
box -33 -37 33 37
use M2M3_PR  M2M3_PR_81
timestamp 1626908933
transform 1 0 240 0 1 14555
box -33 -37 33 37
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_3
timestamp 1626908933
transform 1 0 1700 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_11
timestamp 1626908933
transform 1 0 1700 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_3
timestamp 1626908933
transform 1 0 1700 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_11
timestamp 1626908933
transform 1 0 1700 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_2
timestamp 1626908933
transform 1 0 4100 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_10
timestamp 1626908933
transform 1 0 4100 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_2
timestamp 1626908933
transform 1 0 4100 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_10
timestamp 1626908933
transform 1 0 4100 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA6  prbs_generator_syn_VIA6_0
timestamp 1626908933
transform 1 0 6513 0 1 14636
box -87 -33 87 33
use prbs_generator_syn_VIA6  prbs_generator_syn_VIA6_2
timestamp 1626908933
transform 1 0 6513 0 1 14636
box -87 -33 87 33
use prbs_generator_syn_VIA7  prbs_generator_syn_VIA7_0
timestamp 1626908933
transform 1 0 6513 0 1 14629
box -87 -26 87 26
use prbs_generator_syn_VIA7  prbs_generator_syn_VIA7_2
timestamp 1626908933
transform 1 0 6513 0 1 14629
box -87 -26 87 26
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_1
timestamp 1626908933
transform 1 0 8900 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_9
timestamp 1626908933
transform 1 0 8900 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_1
timestamp 1626908933
transform 1 0 8900 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_9
timestamp 1626908933
transform 1 0 8900 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_0
timestamp 1626908933
transform 1 0 11300 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA4  prbs_generator_syn_VIA4_8
timestamp 1626908933
transform 1 0 11300 0 1 14636
box -100 -33 100 33
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_0
timestamp 1626908933
transform 1 0 11300 0 1 14629
box -100 -26 100 26
use prbs_generator_syn_VIA5  prbs_generator_syn_VIA5_8
timestamp 1626908933
transform 1 0 11300 0 1 14629
box -100 -26 100 26
<< labels >>
rlabel metal2 s 130 0 158 97 4 clk
port 1 nsew
rlabel metal3 s 13856 2691 14016 2751 4 rst
port 2 nsew
rlabel metal3 s 13856 2081 14016 2141 4 cke
port 3 nsew
rlabel metal2 s 898 0 926 97 4 init_val[31]
port 4 nsew
rlabel metal2 s 1666 0 1694 97 4 init_val[30]
port 5 nsew
rlabel metal2 s 2434 0 2462 97 4 init_val[29]
port 6 nsew
rlabel metal2 s 3202 0 3230 97 4 init_val[28]
port 7 nsew
rlabel metal2 s 3970 0 3998 97 4 init_val[27]
port 8 nsew
rlabel metal2 s 4738 0 4766 97 4 init_val[26]
port 9 nsew
rlabel metal2 s 5506 0 5534 97 4 init_val[25]
port 10 nsew
rlabel metal2 s 6274 0 6302 97 4 init_val[24]
port 11 nsew
rlabel metal2 s 7042 0 7070 97 4 init_val[23]
port 12 nsew
rlabel metal2 s 7810 0 7838 97 4 init_val[22]
port 13 nsew
rlabel metal2 s 8578 0 8606 97 4 init_val[21]
port 14 nsew
rlabel metal2 s 9346 0 9374 97 4 init_val[20]
port 15 nsew
rlabel metal2 s 10114 0 10142 97 4 init_val[19]
port 16 nsew
rlabel metal2 s 10882 0 10910 97 4 init_val[18]
port 17 nsew
rlabel metal2 s 11650 0 11678 97 4 init_val[17]
port 18 nsew
rlabel metal2 s 12418 0 12446 97 4 init_val[16]
port 19 nsew
rlabel metal2 s 13186 0 13214 97 4 init_val[15]
port 20 nsew
rlabel metal2 s 13954 0 13982 97 4 init_val[14]
port 21 nsew
rlabel metal3 s 0 14525 160 14585 4 init_val[13]
port 22 nsew
rlabel metal3 s 0 13305 160 13365 4 init_val[12]
port 23 nsew
rlabel metal3 s 0 12207 160 12267 4 init_val[11]
port 24 nsew
rlabel metal3 s 0 11109 160 11169 4 init_val[10]
port 25 nsew
rlabel metal3 s 0 10011 160 10071 4 init_val[9]
port 26 nsew
rlabel metal3 s 0 8913 160 8973 4 init_val[8]
port 27 nsew
rlabel metal3 s 0 7815 160 7875 4 init_val[7]
port 28 nsew
rlabel metal3 s 0 6717 160 6777 4 init_val[6]
port 29 nsew
rlabel metal3 s 0 5619 160 5679 4 init_val[5]
port 30 nsew
rlabel metal3 s 0 4521 160 4581 4 init_val[4]
port 31 nsew
rlabel metal3 s 0 3423 160 3483 4 init_val[3]
port 32 nsew
rlabel metal3 s 0 2325 160 2385 4 init_val[2]
port 33 nsew
rlabel metal3 s 0 1227 160 1287 4 init_val[1]
port 34 nsew
rlabel metal3 s 0 129 160 189 4 init_val[0]
port 35 nsew
rlabel metal3 s 13856 3301 14016 3361 4 eqn[31]
port 36 nsew
rlabel metal3 s 13856 3911 14016 3971 4 eqn[30]
port 37 nsew
rlabel metal3 s 13856 4521 14016 4581 4 eqn[29]
port 38 nsew
rlabel metal3 s 13856 5253 14016 5313 4 eqn[28]
port 39 nsew
rlabel metal3 s 13856 5863 14016 5923 4 eqn[27]
port 40 nsew
rlabel metal3 s 13856 7083 14016 7143 4 eqn[26]
port 41 nsew
rlabel metal3 s 13856 7693 14016 7753 4 eqn[25]
port 42 nsew
rlabel metal3 s 13856 8303 14016 8363 4 eqn[24]
port 43 nsew
rlabel metal3 s 13856 8913 14016 8973 4 eqn[23]
port 44 nsew
rlabel metal3 s 13856 9523 14016 9583 4 eqn[22]
port 45 nsew
rlabel metal3 s 13856 10255 14016 10315 4 eqn[21]
port 46 nsew
rlabel metal3 s 13856 10865 14016 10925 4 eqn[20]
port 47 nsew
rlabel metal3 s 13856 11475 14016 11535 4 eqn[19]
port 48 nsew
rlabel metal3 s 13856 12085 14016 12145 4 eqn[18]
port 49 nsew
rlabel metal3 s 13856 12695 14016 12755 4 eqn[17]
port 50 nsew
rlabel metal3 s 13856 13305 14016 13365 4 eqn[16]
port 51 nsew
rlabel metal3 s 13856 13915 14016 13975 4 eqn[15]
port 52 nsew
rlabel metal3 s 13856 14525 14016 14585 4 eqn[14]
port 53 nsew
rlabel metal2 s 13954 14555 13982 14652 4 eqn[13]
port 54 nsew
rlabel metal2 s 12802 14555 12830 14652 4 eqn[12]
port 55 nsew
rlabel metal2 s 11746 14555 11774 14652 4 eqn[11]
port 56 nsew
rlabel metal2 s 10690 14555 10718 14652 4 eqn[10]
port 57 nsew
rlabel metal2 s 9634 14555 9662 14652 4 eqn[9]
port 58 nsew
rlabel metal2 s 8578 14555 8606 14652 4 eqn[8]
port 59 nsew
rlabel metal2 s 7522 14555 7550 14652 4 eqn[7]
port 60 nsew
rlabel metal2 s 6370 14555 6398 14652 4 eqn[6]
port 61 nsew
rlabel metal2 s 5314 14555 5342 14652 4 eqn[5]
port 62 nsew
rlabel metal2 s 4258 14555 4286 14652 4 eqn[4]
port 63 nsew
rlabel metal2 s 3202 14555 3230 14652 4 eqn[3]
port 64 nsew
rlabel metal2 s 2146 14555 2174 14652 4 eqn[2]
port 65 nsew
rlabel metal2 s 1090 14555 1118 14652 4 eqn[1]
port 66 nsew
rlabel metal2 s 34 14555 62 14652 4 eqn[0]
port 67 nsew
rlabel metal3 s 13856 1471 14016 1531 4 inj_err
port 68 nsew
rlabel metal3 s 13856 251 14016 311 4 inv_chicken[1]
port 69 nsew
rlabel metal3 s 13856 861 14016 921 4 inv_chicken[0]
port 70 nsew
rlabel metal3 s 13856 6473 14016 6533 4 out
port 71 nsew
rlabel metal3 s 1600 0 1800 200 4 DVSS:
port 72 nsew
rlabel metal3 s 1600 14452 1800 14652 4 DVSS:
port 72 nsew
rlabel metal3 s 4000 0 4200 200 4 DVSS:
port 72 nsew
rlabel metal3 s 4000 14452 4200 14652 4 DVSS:
port 72 nsew
rlabel metal3 s 6400 0 6600 200 4 DVSS:
port 72 nsew
rlabel metal3 s 6400 14452 6600 14652 4 DVSS:
port 72 nsew
rlabel metal3 s 8800 0 9000 200 4 DVSS:
port 72 nsew
rlabel metal3 s 8800 14452 9000 14652 4 DVSS:
port 72 nsew
rlabel metal3 s 11200 0 11400 200 4 DVSS:
port 72 nsew
rlabel metal3 s 11200 14452 11400 14652 4 DVSS:
port 72 nsew
rlabel metal1 s 0 -49 98 49 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 -49 14016 49 4 DVSS:
port 72 nsew
rlabel metal1 s 0 1283 98 1381 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 1283 14016 1381 4 DVSS:
port 72 nsew
rlabel metal1 s 0 2615 98 2713 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 2615 14016 2713 4 DVSS:
port 72 nsew
rlabel metal1 s 0 3947 98 4045 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 3947 14016 4045 4 DVSS:
port 72 nsew
rlabel metal1 s 0 5279 98 5377 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 5279 14016 5377 4 DVSS:
port 72 nsew
rlabel metal1 s 0 6611 98 6709 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 6611 14016 6709 4 DVSS:
port 72 nsew
rlabel metal1 s 0 7943 98 8041 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 7943 14016 8041 4 DVSS:
port 72 nsew
rlabel metal1 s 0 9275 98 9373 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 9275 14016 9373 4 DVSS:
port 72 nsew
rlabel metal1 s 0 10607 98 10705 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 10607 14016 10705 4 DVSS:
port 72 nsew
rlabel metal1 s 0 11939 98 12037 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 11939 14016 12037 4 DVSS:
port 72 nsew
rlabel metal1 s 0 13271 98 13369 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 13271 14016 13369 4 DVSS:
port 72 nsew
rlabel metal1 s 0 14603 98 14701 4 DVSS:
port 72 nsew
rlabel metal1 s 13918 14603 14016 14701 4 DVSS:
port 72 nsew
rlabel metal3 s 400 0 600 200 4 DVDD:
port 73 nsew
rlabel metal3 s 400 14452 600 14652 4 DVDD:
port 73 nsew
rlabel metal3 s 2800 0 3000 200 4 DVDD:
port 73 nsew
rlabel metal3 s 2800 14452 3000 14652 4 DVDD:
port 73 nsew
rlabel metal3 s 5200 0 5400 200 4 DVDD:
port 73 nsew
rlabel metal3 s 5200 14452 5400 14652 4 DVDD:
port 73 nsew
rlabel metal3 s 7600 0 7800 200 4 DVDD:
port 73 nsew
rlabel metal3 s 7600 14452 7800 14652 4 DVDD:
port 73 nsew
rlabel metal3 s 10000 0 10200 200 4 DVDD:
port 73 nsew
rlabel metal3 s 10000 14452 10200 14652 4 DVDD:
port 73 nsew
rlabel metal3 s 12400 0 12600 200 4 DVDD:
port 73 nsew
rlabel metal3 s 12400 14452 12600 14652 4 DVDD:
port 73 nsew
rlabel metal1 s 0 617 98 715 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 617 14016 715 4 DVDD:
port 73 nsew
rlabel metal1 s 0 1949 98 2047 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 1949 14016 2047 4 DVDD:
port 73 nsew
rlabel metal1 s 0 3281 98 3379 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 3281 14016 3379 4 DVDD:
port 73 nsew
rlabel metal1 s 0 4613 98 4711 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 4613 14016 4711 4 DVDD:
port 73 nsew
rlabel metal1 s 0 5945 98 6043 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 5945 14016 6043 4 DVDD:
port 73 nsew
rlabel metal1 s 0 7277 98 7375 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 7277 14016 7375 4 DVDD:
port 73 nsew
rlabel metal1 s 0 8609 98 8707 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 8609 14016 8707 4 DVDD:
port 73 nsew
rlabel metal1 s 0 9941 98 10039 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 9941 14016 10039 4 DVDD:
port 73 nsew
rlabel metal1 s 0 11273 98 11371 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 11273 14016 11371 4 DVDD:
port 73 nsew
rlabel metal1 s 0 12605 98 12703 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 12605 14016 12703 4 DVDD:
port 73 nsew
rlabel metal1 s 0 13937 98 14035 4 DVDD:
port 73 nsew
rlabel metal1 s 13918 13937 14016 14035 4 DVDD:
port 73 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 74 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 75 nsew
rlabel metal2 s 144 48 144 48 4 clk
port 1 nsew
rlabel metal3 s 13936 2721 13936 2721 4 rst
port 2 nsew
rlabel metal3 s 13936 2111 13936 2111 4 cke
port 3 nsew
rlabel metal2 s 912 48 912 48 4 init_val[31]
port 4 nsew
rlabel metal2 s 1680 48 1680 48 4 init_val[30]
port 5 nsew
rlabel metal2 s 2448 48 2448 48 4 init_val[29]
port 6 nsew
rlabel metal2 s 3216 48 3216 48 4 init_val[28]
port 7 nsew
rlabel metal2 s 3984 48 3984 48 4 init_val[27]
port 8 nsew
rlabel metal2 s 4752 48 4752 48 4 init_val[26]
port 9 nsew
rlabel metal2 s 5520 48 5520 48 4 init_val[25]
port 10 nsew
rlabel metal2 s 6288 48 6288 48 4 init_val[24]
port 11 nsew
rlabel metal2 s 7056 48 7056 48 4 init_val[23]
port 12 nsew
rlabel metal2 s 7824 48 7824 48 4 init_val[22]
port 13 nsew
rlabel metal2 s 8592 48 8592 48 4 init_val[21]
port 14 nsew
rlabel metal2 s 9360 48 9360 48 4 init_val[20]
port 15 nsew
rlabel metal2 s 10128 48 10128 48 4 init_val[19]
port 16 nsew
rlabel metal2 s 10896 48 10896 48 4 init_val[18]
port 17 nsew
rlabel metal2 s 11664 48 11664 48 4 init_val[17]
port 18 nsew
rlabel metal2 s 12432 48 12432 48 4 init_val[16]
port 19 nsew
rlabel metal2 s 13200 48 13200 48 4 init_val[15]
port 20 nsew
rlabel metal2 s 13968 48 13968 48 4 init_val[14]
port 21 nsew
rlabel metal3 s 80 14555 80 14555 4 init_val[13]
port 22 nsew
rlabel metal3 s 80 13335 80 13335 4 init_val[12]
port 23 nsew
rlabel metal3 s 80 12237 80 12237 4 init_val[11]
port 24 nsew
rlabel metal3 s 80 11139 80 11139 4 init_val[10]
port 25 nsew
rlabel metal3 s 80 10041 80 10041 4 init_val[9]
port 26 nsew
rlabel metal3 s 80 8943 80 8943 4 init_val[8]
port 27 nsew
rlabel metal3 s 80 7845 80 7845 4 init_val[7]
port 28 nsew
rlabel metal3 s 80 6747 80 6747 4 init_val[6]
port 29 nsew
rlabel metal3 s 80 5649 80 5649 4 init_val[5]
port 30 nsew
rlabel metal3 s 80 4551 80 4551 4 init_val[4]
port 31 nsew
rlabel metal3 s 80 3453 80 3453 4 init_val[3]
port 32 nsew
rlabel metal3 s 80 2355 80 2355 4 init_val[2]
port 33 nsew
rlabel metal3 s 80 1257 80 1257 4 init_val[1]
port 34 nsew
rlabel metal3 s 80 159 80 159 4 init_val[0]
port 35 nsew
rlabel metal3 s 13936 3331 13936 3331 4 eqn[31]
port 36 nsew
rlabel metal3 s 13936 3941 13936 3941 4 eqn[30]
port 37 nsew
rlabel metal3 s 13936 4551 13936 4551 4 eqn[29]
port 38 nsew
rlabel metal3 s 13936 5283 13936 5283 4 eqn[28]
port 39 nsew
rlabel metal3 s 13936 5893 13936 5893 4 eqn[27]
port 40 nsew
rlabel metal3 s 13936 7113 13936 7113 4 eqn[26]
port 41 nsew
rlabel metal3 s 13936 7723 13936 7723 4 eqn[25]
port 42 nsew
rlabel metal3 s 13936 8333 13936 8333 4 eqn[24]
port 43 nsew
rlabel metal3 s 13936 8943 13936 8943 4 eqn[23]
port 44 nsew
rlabel metal3 s 13936 9553 13936 9553 4 eqn[22]
port 45 nsew
rlabel metal3 s 13936 10285 13936 10285 4 eqn[21]
port 46 nsew
rlabel metal3 s 13936 10895 13936 10895 4 eqn[20]
port 47 nsew
rlabel metal3 s 13936 11505 13936 11505 4 eqn[19]
port 48 nsew
rlabel metal3 s 13936 12115 13936 12115 4 eqn[18]
port 49 nsew
rlabel metal3 s 13936 12725 13936 12725 4 eqn[17]
port 50 nsew
rlabel metal3 s 13936 13335 13936 13335 4 eqn[16]
port 51 nsew
rlabel metal3 s 13936 13945 13936 13945 4 eqn[15]
port 52 nsew
rlabel metal3 s 13936 14555 13936 14555 4 eqn[14]
port 53 nsew
rlabel metal2 s 13968 14603 13968 14603 4 eqn[13]
port 54 nsew
rlabel metal2 s 12816 14603 12816 14603 4 eqn[12]
port 55 nsew
rlabel metal2 s 11760 14603 11760 14603 4 eqn[11]
port 56 nsew
rlabel metal2 s 10704 14603 10704 14603 4 eqn[10]
port 57 nsew
rlabel metal2 s 9648 14603 9648 14603 4 eqn[9]
port 58 nsew
rlabel metal2 s 8592 14603 8592 14603 4 eqn[8]
port 59 nsew
rlabel metal2 s 7536 14603 7536 14603 4 eqn[7]
port 60 nsew
rlabel metal2 s 6384 14603 6384 14603 4 eqn[6]
port 61 nsew
rlabel metal2 s 5328 14603 5328 14603 4 eqn[5]
port 62 nsew
rlabel metal2 s 4272 14603 4272 14603 4 eqn[4]
port 63 nsew
rlabel metal2 s 3216 14603 3216 14603 4 eqn[3]
port 64 nsew
rlabel metal2 s 2160 14603 2160 14603 4 eqn[2]
port 65 nsew
rlabel metal2 s 1104 14603 1104 14603 4 eqn[1]
port 66 nsew
rlabel metal2 s 48 14603 48 14603 4 eqn[0]
port 67 nsew
rlabel metal3 s 13936 1501 13936 1501 4 inj_err
port 68 nsew
rlabel metal3 s 13936 281 13936 281 4 inv_chicken[1]
port 69 nsew
rlabel metal3 s 13936 891 13936 891 4 inv_chicken[0]
port 70 nsew
rlabel metal3 s 13936 6503 13936 6503 4 out
port 71 nsew
rlabel metal3 s 1700 100 1700 100 4 DVSS:
port 72 nsew
rlabel metal3 s 1700 14552 1700 14552 4 DVSS:
port 72 nsew
rlabel metal3 s 4100 100 4100 100 4 DVSS:
port 72 nsew
rlabel metal3 s 4100 14552 4100 14552 4 DVSS:
port 72 nsew
rlabel metal3 s 6500 100 6500 100 4 DVSS:
port 72 nsew
rlabel metal3 s 6500 14552 6500 14552 4 DVSS:
port 72 nsew
rlabel metal3 s 8900 100 8900 100 4 DVSS:
port 72 nsew
rlabel metal3 s 8900 14552 8900 14552 4 DVSS:
port 72 nsew
rlabel metal3 s 11300 100 11300 100 4 DVSS:
port 72 nsew
rlabel metal3 s 11300 14552 11300 14552 4 DVSS:
port 72 nsew
rlabel metal1 s 49 0 49 0 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 0 13967 0 4 DVSS:
port 72 nsew
rlabel metal1 s 49 1332 49 1332 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 1332 13967 1332 4 DVSS:
port 72 nsew
rlabel metal1 s 49 2664 49 2664 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 2664 13967 2664 4 DVSS:
port 72 nsew
rlabel metal1 s 49 3996 49 3996 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 3996 13967 3996 4 DVSS:
port 72 nsew
rlabel metal1 s 49 5328 49 5328 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 5328 13967 5328 4 DVSS:
port 72 nsew
rlabel metal1 s 49 6660 49 6660 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 6660 13967 6660 4 DVSS:
port 72 nsew
rlabel metal1 s 49 7992 49 7992 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 7992 13967 7992 4 DVSS:
port 72 nsew
rlabel metal1 s 49 9324 49 9324 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 9324 13967 9324 4 DVSS:
port 72 nsew
rlabel metal1 s 49 10656 49 10656 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 10656 13967 10656 4 DVSS:
port 72 nsew
rlabel metal1 s 49 11988 49 11988 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 11988 13967 11988 4 DVSS:
port 72 nsew
rlabel metal1 s 49 13320 49 13320 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 13320 13967 13320 4 DVSS:
port 72 nsew
rlabel metal1 s 49 14652 49 14652 4 DVSS:
port 72 nsew
rlabel metal1 s 13967 14652 13967 14652 4 DVSS:
port 72 nsew
rlabel metal3 s 500 100 500 100 4 DVDD:
port 73 nsew
rlabel metal3 s 500 14552 500 14552 4 DVDD:
port 73 nsew
rlabel metal3 s 2900 100 2900 100 4 DVDD:
port 73 nsew
rlabel metal3 s 2900 14552 2900 14552 4 DVDD:
port 73 nsew
rlabel metal3 s 5300 100 5300 100 4 DVDD:
port 73 nsew
rlabel metal3 s 5300 14552 5300 14552 4 DVDD:
port 73 nsew
rlabel metal3 s 7700 100 7700 100 4 DVDD:
port 73 nsew
rlabel metal3 s 7700 14552 7700 14552 4 DVDD:
port 73 nsew
rlabel metal3 s 10100 100 10100 100 4 DVDD:
port 73 nsew
rlabel metal3 s 10100 14552 10100 14552 4 DVDD:
port 73 nsew
rlabel metal3 s 12500 100 12500 100 4 DVDD:
port 73 nsew
rlabel metal3 s 12500 14552 12500 14552 4 DVDD:
port 73 nsew
rlabel metal1 s 49 666 49 666 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 666 13967 666 4 DVDD:
port 73 nsew
rlabel metal1 s 49 1998 49 1998 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 1998 13967 1998 4 DVDD:
port 73 nsew
rlabel metal1 s 49 3330 49 3330 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 3330 13967 3330 4 DVDD:
port 73 nsew
rlabel metal1 s 49 4662 49 4662 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 4662 13967 4662 4 DVDD:
port 73 nsew
rlabel metal1 s 49 5994 49 5994 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 5994 13967 5994 4 DVDD:
port 73 nsew
rlabel metal1 s 49 7326 49 7326 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 7326 13967 7326 4 DVDD:
port 73 nsew
rlabel metal1 s 49 8658 49 8658 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 8658 13967 8658 4 DVDD:
port 73 nsew
rlabel metal1 s 49 9990 49 9990 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 9990 13967 9990 4 DVDD:
port 73 nsew
rlabel metal1 s 49 11322 49 11322 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 11322 13967 11322 4 DVDD:
port 73 nsew
rlabel metal1 s 49 12654 49 12654 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 12654 13967 12654 4 DVDD:
port 73 nsew
rlabel metal1 s 49 13986 49 13986 4 DVDD:
port 73 nsew
rlabel metal1 s 13967 13986 13967 13986 4 DVDD:
port 73 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 74 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 75 nsew
<< properties >>
string path 140.400 93.425 140.400 97.125 
<< end >>
