magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal2 >>
rect -200 28 200 49
rect -200 -28 -188 28
rect -132 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 132 28
rect 188 -28 200 28
rect -200 -49 200 -28
<< via2 >>
rect -188 -28 -132 28
rect -108 -28 -52 28
rect -28 -28 28 28
rect 52 -28 108 28
rect 132 -28 188 28
<< metal3 >>
rect -200 28 200 49
rect -200 -28 -188 28
rect -132 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 132 28
rect 188 -28 200 28
rect -200 -49 200 -28
<< end >>
