magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 422 704
<< pwell >>
rect 0 0 384 49
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 0 617 384 666 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 0 0 384 49 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
flabel pwell s 192 24 192 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 192 641 192 641 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 fill_4
flabel metal1 s 192 641 192 641 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 192 24 192 24 0 FreeSans 200 0 0 0 VGND
<< properties >>
string FIXED_BBOX 0 0 384 666
<< end >>
