magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal3 >>
rect -200 32 200 33
rect -200 -32 -192 32
rect -128 -32 -112 32
rect -48 -32 -32 32
rect 32 -32 48 32
rect 112 -32 128 32
rect 192 -32 200 32
rect -200 -33 200 -32
<< via3 >>
rect -192 -32 -128 32
rect -112 -32 -48 32
rect -32 -32 32 32
rect 48 -32 112 32
rect 128 -32 192 32
<< metal4 >>
rect -200 32 200 33
rect -200 -32 -192 32
rect -128 -32 -112 32
rect -48 -32 -32 32
rect 32 -32 48 32
rect 112 -32 128 32
rect 192 -32 200 32
rect -200 -33 200 -32
<< end >>
