magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal2 >>
rect -292 28 292 49
rect -292 -28 -268 28
rect -212 -28 -188 28
rect -132 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 132 28
rect 188 -28 212 28
rect 268 -28 292 28
rect -292 -49 292 -28
<< via2 >>
rect -268 -28 -212 28
rect -188 -28 -132 28
rect -108 -28 -52 28
rect -28 -28 28 28
rect 52 -28 108 28
rect 132 -28 188 28
rect 212 -28 268 28
<< metal3 >>
rect -292 28 292 49
rect -292 -28 -268 28
rect -212 -28 -188 28
rect -132 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 132 28
rect 188 -28 212 28
rect 268 -28 292 28
rect -292 -49 292 -28
<< end >>
