magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 0 0 960 49
<< scpmos >>
rect 87 368 117 592
rect 185 368 215 592
rect 283 368 313 592
rect 377 368 407 592
rect 539 368 569 592
rect 629 368 659 592
rect 741 368 771 592
rect 831 368 861 592
<< nmoslvt >>
rect 84 74 114 222
rect 188 74 218 222
rect 274 74 304 222
rect 360 74 390 222
rect 572 74 602 222
rect 658 74 688 222
rect 744 74 774 222
rect 834 74 864 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 144 188 222
rect 114 110 139 144
rect 173 110 188 144
rect 114 74 188 110
rect 218 210 274 222
rect 218 176 229 210
rect 263 176 274 210
rect 218 120 274 176
rect 218 86 229 120
rect 263 86 274 120
rect 218 74 274 86
rect 304 189 360 222
rect 304 155 315 189
rect 349 155 360 189
rect 304 74 360 155
rect 390 164 440 222
rect 390 136 461 164
rect 522 150 572 222
rect 390 102 415 136
rect 449 102 461 136
rect 390 74 461 102
rect 515 142 572 150
rect 515 108 527 142
rect 561 108 572 142
rect 515 74 572 108
rect 602 179 658 222
rect 602 145 613 179
rect 647 145 658 179
rect 602 74 658 145
rect 688 210 744 222
rect 688 176 699 210
rect 733 176 744 210
rect 688 120 744 176
rect 688 86 699 120
rect 733 86 744 120
rect 688 74 744 86
rect 774 179 834 222
rect 774 145 785 179
rect 819 145 834 179
rect 774 74 834 145
rect 864 164 914 222
rect 864 136 931 164
rect 864 102 885 136
rect 919 102 931 136
rect 864 74 931 102
<< pdiff >>
rect 27 580 87 592
rect 27 546 39 580
rect 73 546 87 580
rect 27 503 87 546
rect 27 469 39 503
rect 73 469 87 503
rect 27 424 87 469
rect 27 390 39 424
rect 73 390 87 424
rect 27 368 87 390
rect 117 580 185 592
rect 117 546 130 580
rect 164 546 185 580
rect 117 508 185 546
rect 117 474 130 508
rect 164 474 185 508
rect 117 440 185 474
rect 117 406 130 440
rect 164 406 185 440
rect 117 368 185 406
rect 215 580 283 592
rect 215 546 230 580
rect 264 546 283 580
rect 215 499 283 546
rect 215 465 230 499
rect 264 465 283 499
rect 215 368 283 465
rect 313 580 377 592
rect 313 546 330 580
rect 364 546 377 580
rect 313 503 377 546
rect 313 469 330 503
rect 364 469 377 503
rect 313 424 377 469
rect 313 390 330 424
rect 364 390 377 424
rect 313 368 377 390
rect 407 580 539 592
rect 407 546 420 580
rect 454 546 492 580
rect 526 546 539 580
rect 407 508 539 546
rect 407 474 420 508
rect 454 474 492 508
rect 526 474 539 508
rect 407 368 539 474
rect 569 580 629 592
rect 569 546 582 580
rect 616 546 629 580
rect 569 503 629 546
rect 569 469 582 503
rect 616 469 629 503
rect 569 424 629 469
rect 569 390 582 424
rect 616 390 629 424
rect 569 368 629 390
rect 659 580 741 592
rect 659 546 682 580
rect 716 546 741 580
rect 659 499 741 546
rect 659 465 682 499
rect 716 465 741 499
rect 659 368 741 465
rect 771 580 831 592
rect 771 546 784 580
rect 818 546 831 580
rect 771 503 831 546
rect 771 469 784 503
rect 818 469 831 503
rect 771 424 831 469
rect 771 390 784 424
rect 818 390 831 424
rect 771 368 831 390
rect 861 580 924 592
rect 861 546 875 580
rect 909 546 924 580
rect 861 499 924 546
rect 861 465 875 499
rect 909 465 924 499
rect 861 368 924 465
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 110 173 144
rect 229 176 263 210
rect 229 86 263 120
rect 315 155 349 189
rect 415 102 449 136
rect 527 108 561 142
rect 613 145 647 179
rect 699 176 733 210
rect 699 86 733 120
rect 785 145 819 179
rect 885 102 919 136
<< pdiffc >>
rect 39 546 73 580
rect 39 469 73 503
rect 39 390 73 424
rect 130 546 164 580
rect 130 474 164 508
rect 130 406 164 440
rect 230 546 264 580
rect 230 465 264 499
rect 330 546 364 580
rect 330 469 364 503
rect 330 390 364 424
rect 420 546 454 580
rect 492 546 526 580
rect 420 474 454 508
rect 492 474 526 508
rect 582 546 616 580
rect 582 469 616 503
rect 582 390 616 424
rect 682 546 716 580
rect 682 465 716 499
rect 784 546 818 580
rect 784 469 818 503
rect 784 390 818 424
rect 875 546 909 580
rect 875 465 909 499
<< poly >>
rect 87 592 117 618
rect 185 592 215 618
rect 283 592 313 618
rect 377 592 407 618
rect 539 592 569 618
rect 629 592 659 618
rect 741 592 771 618
rect 831 592 861 618
rect 87 353 117 368
rect 185 353 215 368
rect 283 353 313 368
rect 377 353 407 368
rect 539 353 569 368
rect 629 353 659 368
rect 741 353 771 368
rect 831 353 861 368
rect 84 336 120 353
rect 182 336 218 353
rect 84 320 218 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 218 320
rect 280 336 316 353
rect 374 336 410 353
rect 536 336 572 353
rect 626 336 662 353
rect 741 336 774 353
rect 828 336 864 353
rect 280 320 488 336
rect 280 300 302 320
rect 84 270 218 286
rect 84 222 114 270
rect 188 222 218 270
rect 274 286 302 300
rect 336 286 370 320
rect 404 286 438 320
rect 472 286 488 320
rect 274 270 488 286
rect 536 320 688 336
rect 536 286 552 320
rect 586 286 638 320
rect 672 286 688 320
rect 536 270 688 286
rect 274 222 304 270
rect 360 222 390 270
rect 572 222 602 270
rect 658 222 688 270
rect 744 320 864 336
rect 744 286 793 320
rect 827 286 864 320
rect 744 270 864 286
rect 744 222 774 270
rect 834 222 864 270
rect 84 48 114 74
rect 188 48 218 74
rect 274 48 304 74
rect 360 48 390 74
rect 572 48 602 74
rect 658 48 688 74
rect 744 48 774 74
rect 834 48 864 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 302 286 336 320
rect 370 286 404 320
rect 438 286 472 320
rect 552 286 586 320
rect 638 286 672 320
rect 793 286 827 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 90 649
rect 23 546 39 580
rect 73 546 90 580
rect 23 503 90 546
rect 23 469 39 503
rect 73 469 90 503
rect 23 424 90 469
rect 23 390 39 424
rect 73 390 90 424
rect 127 580 180 596
rect 127 546 130 580
rect 164 546 180 580
rect 127 508 180 546
rect 127 474 130 508
rect 164 474 180 508
rect 127 440 180 474
rect 214 580 280 649
rect 214 546 230 580
rect 264 546 280 580
rect 214 499 280 546
rect 214 465 230 499
rect 264 465 280 499
rect 214 458 280 465
rect 314 580 380 596
rect 314 546 330 580
rect 364 546 380 580
rect 314 503 380 546
rect 314 469 330 503
rect 364 469 380 503
rect 127 406 130 440
rect 164 424 180 440
rect 314 424 380 469
rect 416 580 530 649
rect 416 546 420 580
rect 454 546 492 580
rect 526 546 530 580
rect 416 508 530 546
rect 416 474 420 508
rect 454 474 492 508
rect 526 474 530 508
rect 416 458 530 474
rect 566 580 632 596
rect 566 546 582 580
rect 616 546 632 580
rect 566 503 632 546
rect 566 469 582 503
rect 616 469 632 503
rect 566 424 632 469
rect 666 580 732 649
rect 666 546 682 580
rect 716 546 732 580
rect 666 499 732 546
rect 666 465 682 499
rect 716 465 732 499
rect 666 458 732 465
rect 768 580 825 596
rect 768 546 784 580
rect 818 546 825 580
rect 768 503 825 546
rect 768 469 784 503
rect 818 469 825 503
rect 768 430 825 469
rect 859 580 925 649
rect 859 546 875 580
rect 909 546 925 580
rect 859 499 925 546
rect 859 465 875 499
rect 909 465 925 499
rect 859 464 925 465
rect 768 424 935 430
rect 164 406 330 424
rect 127 390 330 406
rect 364 390 582 424
rect 616 390 784 424
rect 818 390 935 424
rect 25 320 218 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 218 320
rect 25 270 218 286
rect 286 320 488 356
rect 286 286 302 320
rect 336 286 370 320
rect 404 286 438 320
rect 472 286 488 320
rect 286 270 488 286
rect 536 320 743 356
rect 536 286 552 320
rect 586 286 638 320
rect 672 286 743 320
rect 536 270 743 286
rect 777 320 843 356
rect 777 286 793 320
rect 827 286 843 320
rect 777 270 843 286
rect 889 236 935 390
rect 23 210 263 236
rect 23 176 39 210
rect 73 202 229 210
rect 73 176 89 202
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 144 189 168
rect 123 110 139 144
rect 173 110 189 144
rect 123 17 189 110
rect 229 120 263 176
rect 299 202 663 236
rect 299 189 365 202
rect 299 155 315 189
rect 349 155 365 189
rect 597 179 663 202
rect 299 119 365 155
rect 399 136 465 168
rect 229 85 263 86
rect 399 102 415 136
rect 449 102 465 136
rect 399 85 465 102
rect 229 51 465 85
rect 511 142 563 168
rect 511 108 527 142
rect 561 108 563 142
rect 597 145 613 179
rect 647 145 663 179
rect 597 129 663 145
rect 697 210 735 226
rect 697 176 699 210
rect 733 176 735 210
rect 511 85 563 108
rect 697 120 735 176
rect 769 202 935 236
rect 769 179 835 202
rect 769 145 785 179
rect 819 145 835 179
rect 769 129 835 145
rect 869 136 935 168
rect 697 86 699 120
rect 733 86 735 120
rect 697 85 735 86
rect 869 102 885 136
rect 919 102 935 136
rect 869 85 935 102
rect 511 51 935 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4_2
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
rlabel comment s 0 0 0 0 4 nand4_2
flabel pwell s 480 24 480 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 480 641 480 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 480 641 480 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 480 24 480 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 912 259 912 259 0 FreeSans 340 0 0 0 Y
flabel locali s 912 333 912 333 0 FreeSans 340 0 0 0 Y
flabel locali s 912 407 912 407 0 FreeSans 340 0 0 0 Y
flabel locali s 336 333 336 333 0 FreeSans 340 0 0 0 C
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 C
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 D
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 D
flabel locali s 624 333 624 333 0 FreeSans 340 0 0 0 B
flabel locali s 720 333 720 333 0 FreeSans 340 0 0 0 B
flabel locali s 816 333 816 333 0 FreeSans 340 0 0 0 A
rlabel comment s 0 0 0 0 4 nand4_2
flabel pwell s 480 24 480 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 480 641 480 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 480 641 480 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 480 24 480 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 912 259 912 259 0 FreeSans 340 0 0 0 Y
flabel locali s 912 333 912 333 0 FreeSans 340 0 0 0 Y
flabel locali s 912 407 912 407 0 FreeSans 340 0 0 0 Y
flabel locali s 336 333 336 333 0 FreeSans 340 0 0 0 C
flabel locali s 432 333 432 333 0 FreeSans 340 0 0 0 C
flabel locali s 48 333 48 333 0 FreeSans 340 0 0 0 D
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 D
flabel locali s 624 333 624 333 0 FreeSans 340 0 0 0 B
flabel locali s 720 333 720 333 0 FreeSans 340 0 0 0 B
flabel locali s 816 333 816 333 0 FreeSans 340 0 0 0 A
<< properties >>
string FIXED_BBOX 0 0 960 666
<< end >>
