magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< error_s >>
rect 1118 19835 1119 19880
rect 2078 19835 2079 19880
rect 5630 19835 5631 19880
rect 8894 19835 8895 19880
rect 10142 19835 10143 19880
rect 11390 19835 11391 19880
rect 14654 19835 14655 19880
rect 15902 19835 15903 19880
rect 16958 19835 16959 19880
rect 19166 19835 19167 19880
rect 20414 19835 20415 19880
rect 23006 19835 23007 19880
rect 24254 19835 24255 19880
rect 25598 19835 25599 19880
rect 26846 19835 26847 19880
rect 28190 19835 28191 19880
rect 29438 19835 29439 19880
rect 30686 19835 30687 19880
rect 32030 19835 32031 19880
rect 33278 19835 33279 19880
rect 34526 19835 34527 19880
rect 35294 19835 35295 19880
rect 10814 18759 10815 18804
rect 15614 18759 15615 18804
rect 24254 18759 24255 18804
rect 25598 18759 25599 18804
rect 26846 18759 26847 18804
rect 28190 18759 28191 18804
rect 29438 18759 29439 18804
rect 30686 18759 30687 18804
rect 32030 18759 32031 18804
rect 33278 18759 33279 18804
rect 34526 18759 34527 18804
rect 638 18503 639 18548
rect 10814 18503 10815 18548
rect 15614 18503 15615 18548
rect 19742 18503 19743 18548
rect 23678 18503 23679 18548
rect 24926 18503 24927 18548
rect 26174 18503 26175 18548
rect 27038 18503 27039 18548
rect 28190 18503 28191 18548
rect 29438 18503 29439 18548
rect 30686 18503 30687 18548
rect 32030 18503 32031 18548
rect 33278 18503 33279 18548
rect 34526 18503 34527 18548
rect 35294 18503 35295 18548
rect 2462 17427 2463 17472
rect 6974 17427 6975 17472
rect 8606 17427 8607 17472
rect 10814 17427 10815 17472
rect 12734 17427 12735 17472
rect 14558 17427 14559 17472
rect 15614 17427 15615 17472
rect 17246 17427 17247 17472
rect 19166 17427 19167 17472
rect 21566 17427 21567 17472
rect 23678 17427 23679 17472
rect 24542 17427 24543 17472
rect 25598 17427 25599 17472
rect 26846 17427 26847 17472
rect 28190 17427 28191 17472
rect 29438 17427 29439 17472
rect 30686 17427 30687 17472
rect 32030 17427 32031 17472
rect 33278 17427 33279 17472
rect 34526 17427 34527 17472
rect 638 17171 639 17216
rect 2078 17171 2079 17216
rect 6974 17171 6975 17216
rect 15326 17171 15327 17216
rect 17054 17171 17055 17216
rect 19166 17171 19167 17216
rect 21086 17171 21087 17216
rect 23006 17171 23007 17216
rect 24254 17171 24255 17216
rect 25598 17171 25599 17216
rect 26846 17171 26847 17216
rect 28190 17171 28191 17216
rect 29438 17171 29439 17216
rect 30686 17171 30687 17216
rect 32030 17171 32031 17216
rect 33278 17171 33279 17216
rect 34526 17171 34527 17216
rect 35294 17171 35295 17216
rect 2462 16095 2463 16140
rect 4574 16095 4575 16140
rect 10814 16095 10815 16140
rect 12734 16095 12735 16140
rect 13982 16095 13983 16140
rect 15614 16095 15615 16140
rect 17054 16095 17055 16140
rect 19166 16095 19167 16140
rect 21086 16095 21087 16140
rect 23006 16095 23007 16140
rect 25598 16095 25599 16140
rect 26846 16095 26847 16140
rect 28190 16095 28191 16140
rect 29438 16095 29439 16140
rect 30686 16095 30687 16140
rect 32030 16095 32031 16140
rect 33278 16095 33279 16140
rect 34526 16095 34527 16140
rect 15326 15839 15327 15884
rect 16574 15839 16575 15884
rect 19742 15839 19743 15884
rect 20990 15839 20991 15884
rect 23678 15839 23679 15884
rect 26174 15839 26175 15884
rect 26942 15839 26943 15884
rect 30686 15839 30687 15884
rect 32030 15839 32031 15884
rect 33278 15839 33279 15884
rect 34526 15839 34527 15884
rect 35294 15839 35295 15884
rect 7166 14763 7167 14808
rect 15902 14763 15903 14808
rect 17054 14763 17055 14808
rect 19550 14763 19551 14808
rect 20414 14763 20415 14808
rect 23616 14785 23617 14796
rect 25728 14785 25729 14796
rect 23627 14751 23628 14785
rect 25739 14751 25740 14785
rect 30686 14763 30687 14808
rect 32030 14763 32031 14808
rect 33278 14763 33279 14808
rect 34526 14763 34527 14808
rect 23424 14553 23425 14564
rect 15326 14507 15327 14552
rect 16574 14507 16575 14552
rect 19742 14507 19743 14552
rect 20990 14507 20991 14552
rect 23435 14519 23436 14553
rect 30686 14507 30687 14552
rect 32030 14507 32031 14552
rect 33278 14507 33279 14552
rect 34526 14507 34527 14552
rect 35294 14507 35295 14552
rect 15902 13431 15903 13476
rect 17054 13431 17055 13476
rect 19550 13431 19551 13476
rect 20414 13431 20415 13476
rect 32030 13431 32031 13476
rect 33278 13431 33279 13476
rect 34526 13431 34527 13476
rect 26208 13221 26209 13232
rect 26976 13221 26977 13232
rect 15326 13175 15327 13220
rect 16574 13175 16575 13220
rect 19742 13175 19743 13220
rect 20990 13175 20991 13220
rect 26219 13187 26220 13221
rect 26987 13187 26988 13221
rect 28190 13175 28191 13220
rect 29246 13175 29247 13220
rect 32030 13175 32031 13220
rect 33278 13175 33279 13220
rect 34526 13175 34527 13220
rect 35294 13175 35295 13220
rect 13310 12099 13311 12144
rect 15902 12099 15903 12144
rect 17054 12099 17055 12144
rect 18494 12099 18495 12144
rect 19550 12099 19551 12144
rect 20414 12099 20415 12144
rect 21758 12099 21759 12144
rect 22848 12121 22849 12132
rect 23616 12121 23617 12132
rect 26400 12121 26401 12132
rect 22859 12087 22860 12121
rect 23627 12087 23628 12121
rect 26411 12087 26412 12121
rect 32030 12099 32031 12144
rect 33278 12099 33279 12144
rect 34526 12099 34527 12144
rect 22944 11889 22945 11900
rect 23712 11889 23713 11900
rect 26496 11889 26497 11900
rect 15902 11843 15903 11888
rect 17054 11843 17055 11888
rect 18494 11843 18495 11888
rect 19742 11843 19743 11888
rect 21086 11843 21087 11888
rect 22046 11843 22047 11888
rect 22955 11855 22956 11889
rect 23723 11855 23724 11889
rect 26507 11855 26508 11889
rect 28190 11843 28191 11888
rect 29246 11843 29247 11888
rect 32030 11843 32031 11888
rect 33278 11843 33279 11888
rect 34526 11843 34527 11888
rect 35294 11843 35295 11888
rect 5534 10767 5535 10812
rect 8222 10767 8223 10812
rect 11390 10767 11391 10812
rect 15902 10767 15903 10812
rect 17246 10767 17247 10812
rect 18494 10767 18495 10812
rect 19550 10767 19551 10812
rect 20414 10767 20415 10812
rect 21758 10767 21759 10812
rect 22910 10767 22911 10812
rect 23616 10789 23617 10800
rect 26592 10789 26593 10800
rect 23627 10755 23628 10789
rect 26603 10755 26604 10789
rect 28766 10767 28767 10812
rect 32030 10767 32031 10812
rect 33278 10767 33279 10812
rect 34526 10767 34527 10812
rect 9278 10511 9279 10556
rect 14654 10511 14655 10556
rect 15902 10511 15903 10556
rect 17054 10511 17055 10556
rect 18494 10511 18495 10556
rect 19742 10511 19743 10556
rect 21086 10511 21087 10556
rect 22046 10511 22047 10556
rect 23006 10511 23007 10556
rect 23774 10511 23775 10556
rect 29918 10511 29919 10556
rect 31358 10511 31359 10556
rect 33278 10511 33279 10556
rect 34526 10511 34527 10556
rect 35294 10511 35295 10556
rect 1790 9435 1791 9480
rect 2558 9435 2559 9480
rect 5438 9435 5439 9480
rect 10526 9435 10527 9480
rect 12734 9435 12735 9480
rect 13982 9435 13983 9480
rect 15902 9435 15903 9480
rect 17246 9435 17247 9480
rect 18494 9435 18495 9480
rect 19550 9435 19551 9480
rect 20414 9435 20415 9480
rect 21758 9435 21759 9480
rect 23006 9435 23007 9480
rect 24254 9435 24255 9480
rect 25598 9435 25599 9480
rect 26846 9435 26847 9480
rect 28190 9435 28191 9480
rect 29438 9435 29439 9480
rect 30686 9435 30687 9480
rect 32030 9435 32031 9480
rect 33278 9435 33279 9480
rect 34526 9435 34527 9480
rect 1790 9179 1791 9224
rect 11390 9179 11391 9224
rect 13310 9179 13311 9224
rect 14654 9179 14655 9224
rect 15902 9179 15903 9224
rect 17054 9179 17055 9224
rect 18494 9179 18495 9224
rect 19742 9179 19743 9224
rect 21086 9179 21087 9224
rect 22046 9179 22047 9224
rect 23006 9179 23007 9224
rect 24254 9179 24255 9224
rect 25598 9179 25599 9224
rect 26846 9179 26847 9224
rect 28190 9179 28191 9224
rect 29438 9179 29439 9224
rect 30686 9179 30687 9224
rect 32030 9179 32031 9224
rect 33278 9179 33279 9224
rect 34526 9179 34527 9224
rect 35294 9179 35295 9224
rect 1502 8103 1503 8148
rect 4382 8103 4383 8148
rect 6974 8103 6975 8148
rect 10814 8103 10815 8148
rect 12062 8103 12063 8148
rect 13310 8103 13311 8148
rect 14558 8103 14559 8148
rect 15902 8103 15903 8148
rect 17246 8103 17247 8148
rect 18494 8103 18495 8148
rect 19550 8103 19551 8148
rect 20414 8103 20415 8148
rect 21758 8103 21759 8148
rect 23006 8103 23007 8148
rect 24254 8103 24255 8148
rect 25598 8103 25599 8148
rect 26846 8103 26847 8148
rect 28190 8103 28191 8148
rect 29438 8103 29439 8148
rect 30686 8103 30687 8148
rect 32030 8103 32031 8148
rect 33278 8103 33279 8148
rect 34526 8103 34527 8148
rect 1790 7847 1791 7892
rect 4382 7847 4383 7892
rect 5342 7847 5343 7892
rect 6974 7847 6975 7892
rect 10142 7847 10143 7892
rect 11390 7847 11391 7892
rect 13310 7847 13311 7892
rect 14654 7847 14655 7892
rect 15902 7847 15903 7892
rect 17054 7847 17055 7892
rect 18494 7847 18495 7892
rect 19742 7847 19743 7892
rect 21086 7847 21087 7892
rect 22046 7847 22047 7892
rect 23006 7847 23007 7892
rect 24254 7847 24255 7892
rect 25598 7847 25599 7892
rect 26846 7847 26847 7892
rect 28190 7847 28191 7892
rect 29438 7847 29439 7892
rect 30686 7847 30687 7892
rect 32030 7847 32031 7892
rect 33278 7847 33279 7892
rect 34526 7847 34527 7892
rect 35294 7847 35295 7892
rect 2462 6771 2463 6816
rect 4382 6771 4383 6816
rect 6974 6771 6975 6816
rect 8222 6771 8223 6816
rect 10814 6771 10815 6816
rect 12062 6771 12063 6816
rect 13310 6771 13311 6816
rect 14558 6771 14559 6816
rect 15902 6771 15903 6816
rect 17246 6771 17247 6816
rect 18494 6771 18495 6816
rect 19550 6771 19551 6816
rect 20414 6771 20415 6816
rect 21758 6771 21759 6816
rect 23006 6771 23007 6816
rect 24254 6771 24255 6816
rect 25598 6771 25599 6816
rect 26846 6771 26847 6816
rect 28190 6771 28191 6816
rect 29438 6771 29439 6816
rect 30686 6771 30687 6816
rect 32030 6771 32031 6816
rect 33278 6771 33279 6816
rect 34526 6771 34527 6816
rect 1790 6515 1791 6560
rect 4382 6515 4383 6560
rect 5630 6515 5631 6560
rect 6974 6515 6975 6560
rect 8222 6515 8223 6560
rect 9470 6515 9471 6560
rect 10814 6515 10815 6560
rect 12062 6515 12063 6560
rect 13310 6515 13311 6560
rect 14654 6515 14655 6560
rect 15902 6515 15903 6560
rect 17054 6515 17055 6560
rect 18494 6515 18495 6560
rect 19742 6515 19743 6560
rect 21086 6515 21087 6560
rect 22046 6515 22047 6560
rect 23006 6515 23007 6560
rect 24254 6515 24255 6560
rect 25598 6515 25599 6560
rect 26846 6515 26847 6560
rect 28190 6515 28191 6560
rect 29438 6515 29439 6560
rect 30686 6515 30687 6560
rect 32030 6515 32031 6560
rect 33278 6515 33279 6560
rect 34526 6515 34527 6560
rect 35294 6515 35295 6560
rect 1790 5439 1791 5484
rect 2558 5439 2559 5484
rect 4382 5439 4383 5484
rect 5630 5439 5631 5484
rect 6974 5439 6975 5484
rect 8222 5439 8223 5484
rect 9470 5439 9471 5484
rect 10814 5439 10815 5484
rect 12062 5439 12063 5484
rect 13310 5439 13311 5484
rect 14558 5439 14559 5484
rect 15902 5439 15903 5484
rect 17246 5439 17247 5484
rect 18494 5439 18495 5484
rect 19550 5439 19551 5484
rect 20414 5439 20415 5484
rect 21758 5439 21759 5484
rect 23006 5439 23007 5484
rect 24254 5439 24255 5484
rect 25598 5439 25599 5484
rect 26846 5439 26847 5484
rect 28190 5439 28191 5484
rect 29438 5439 29439 5484
rect 30686 5439 30687 5484
rect 32030 5439 32031 5484
rect 33278 5439 33279 5484
rect 34526 5439 34527 5484
rect 1790 5183 1791 5228
rect 3038 5183 3039 5228
rect 4382 5183 4383 5228
rect 5630 5183 5631 5228
rect 6974 5183 6975 5228
rect 8222 5183 8223 5228
rect 9470 5183 9471 5228
rect 10814 5183 10815 5228
rect 12062 5183 12063 5228
rect 13310 5183 13311 5228
rect 14654 5183 14655 5228
rect 15902 5183 15903 5228
rect 17054 5183 17055 5228
rect 18494 5183 18495 5228
rect 19742 5183 19743 5228
rect 21086 5183 21087 5228
rect 22046 5183 22047 5228
rect 23006 5183 23007 5228
rect 24254 5183 24255 5228
rect 25598 5183 25599 5228
rect 26846 5183 26847 5228
rect 28190 5183 28191 5228
rect 29438 5183 29439 5228
rect 30686 5183 30687 5228
rect 32030 5183 32031 5228
rect 33278 5183 33279 5228
rect 34526 5183 34527 5228
rect 35294 5183 35295 5228
rect 1790 4107 1791 4152
rect 3038 4107 3039 4152
rect 4382 4107 4383 4152
rect 5630 4107 5631 4152
rect 6974 4107 6975 4152
rect 8222 4107 8223 4152
rect 9470 4107 9471 4152
rect 10814 4107 10815 4152
rect 12062 4107 12063 4152
rect 13310 4107 13311 4152
rect 14558 4107 14559 4152
rect 15902 4107 15903 4152
rect 17246 4107 17247 4152
rect 18494 4107 18495 4152
rect 19550 4107 19551 4152
rect 20414 4107 20415 4152
rect 21758 4107 21759 4152
rect 23006 4107 23007 4152
rect 24254 4107 24255 4152
rect 25598 4107 25599 4152
rect 26846 4107 26847 4152
rect 28190 4107 28191 4152
rect 29438 4107 29439 4152
rect 30686 4107 30687 4152
rect 32030 4107 32031 4152
rect 33278 4107 33279 4152
rect 34526 4107 34527 4152
rect 734 3851 735 3896
rect 2078 3851 2079 3896
rect 3038 3851 3039 3896
rect 4382 3851 4383 3896
rect 5630 3851 5631 3896
rect 6974 3851 6975 3896
rect 8222 3851 8223 3896
rect 9470 3851 9471 3896
rect 10814 3851 10815 3896
rect 12062 3851 12063 3896
rect 13310 3851 13311 3896
rect 14654 3851 14655 3896
rect 15902 3851 15903 3896
rect 17054 3851 17055 3896
rect 18494 3851 18495 3896
rect 19742 3851 19743 3896
rect 21086 3851 21087 3896
rect 22046 3851 22047 3896
rect 23006 3851 23007 3896
rect 24254 3851 24255 3896
rect 25598 3851 25599 3896
rect 26846 3851 26847 3896
rect 28190 3851 28191 3896
rect 29438 3851 29439 3896
rect 30686 3851 30687 3896
rect 32030 3851 32031 3896
rect 33278 3851 33279 3896
rect 34526 3851 34527 3896
rect 35294 3851 35295 3896
rect 672 2797 673 2808
rect 683 2763 684 2797
rect 3038 2775 3039 2820
rect 4382 2775 4383 2820
rect 5630 2775 5631 2820
rect 6974 2775 6975 2820
rect 8222 2775 8223 2820
rect 9470 2775 9471 2820
rect 10814 2775 10815 2820
rect 12062 2775 12063 2820
rect 13310 2775 13311 2820
rect 14558 2775 14559 2820
rect 15902 2775 15903 2820
rect 17246 2775 17247 2820
rect 18494 2775 18495 2820
rect 19550 2775 19551 2820
rect 20414 2775 20415 2820
rect 21758 2775 21759 2820
rect 23006 2775 23007 2820
rect 24254 2775 24255 2820
rect 25598 2775 25599 2820
rect 26846 2775 26847 2820
rect 28190 2775 28191 2820
rect 29438 2775 29439 2820
rect 30686 2775 30687 2820
rect 32030 2775 32031 2820
rect 33278 2775 33279 2820
rect 34526 2775 34527 2820
rect 672 2565 673 2576
rect 1440 2565 1441 2576
rect 16992 2565 16993 2576
rect 683 2531 684 2565
rect 1451 2531 1452 2565
rect 3710 2519 3711 2564
rect 4958 2519 4959 2564
rect 6302 2519 6303 2564
rect 7070 2519 7071 2564
rect 8222 2519 8223 2564
rect 9470 2519 9471 2564
rect 10814 2519 10815 2564
rect 12062 2519 12063 2564
rect 13310 2519 13311 2564
rect 14654 2519 14655 2564
rect 15902 2519 15903 2564
rect 17003 2531 17004 2565
rect 18494 2519 18495 2564
rect 19742 2519 19743 2564
rect 21086 2519 21087 2564
rect 22046 2519 22047 2564
rect 23006 2519 23007 2564
rect 24254 2519 24255 2564
rect 25598 2519 25599 2564
rect 26846 2519 26847 2564
rect 28190 2519 28191 2564
rect 29438 2519 29439 2564
rect 30686 2519 30687 2564
rect 32030 2519 32031 2564
rect 33278 2519 33279 2564
rect 34526 2519 34527 2564
rect 35294 2519 35295 2564
rect 672 1465 673 1476
rect 1440 1465 1441 1476
rect 2208 1465 2209 1476
rect 683 1431 684 1465
rect 1451 1431 1452 1465
rect 2219 1431 2220 1465
rect 4382 1443 4383 1488
rect 5630 1443 5631 1488
rect 6974 1443 6975 1488
rect 8222 1443 8223 1488
rect 9470 1443 9471 1488
rect 10814 1443 10815 1488
rect 12062 1443 12063 1488
rect 13310 1443 13311 1488
rect 15710 1443 15711 1488
rect 16416 1465 16417 1476
rect 17184 1465 17185 1476
rect 17952 1465 17953 1476
rect 16427 1431 16428 1465
rect 17195 1431 17196 1465
rect 17963 1431 17964 1465
rect 19166 1443 19167 1488
rect 20414 1443 20415 1488
rect 21758 1443 21759 1488
rect 23006 1443 23007 1488
rect 24254 1443 24255 1488
rect 25598 1443 25599 1488
rect 26846 1443 26847 1488
rect 28190 1443 28191 1488
rect 29438 1443 29439 1488
rect 30686 1443 30687 1488
rect 32030 1443 32031 1488
rect 33278 1443 33279 1488
rect 34526 1443 34527 1488
rect 576 1233 577 1244
rect 1440 1233 1441 1244
rect 13344 1233 13345 1244
rect 14112 1233 14113 1244
rect 14880 1233 14881 1244
rect 15648 1233 15649 1244
rect 16416 1233 16417 1244
rect 17952 1233 17953 1244
rect 587 1199 588 1233
rect 1451 1199 1452 1233
rect 4958 1187 4959 1232
rect 6302 1187 6303 1232
rect 7070 1187 7071 1232
rect 8222 1187 8223 1232
rect 9470 1187 9471 1232
rect 10814 1187 10815 1232
rect 12062 1187 12063 1232
rect 13355 1199 13356 1233
rect 14123 1199 14124 1233
rect 14891 1199 14892 1233
rect 15659 1199 15660 1233
rect 16427 1199 16428 1233
rect 17963 1199 17964 1233
rect 19166 1187 19167 1232
rect 20414 1187 20415 1232
rect 21758 1187 21759 1232
rect 23006 1187 23007 1232
rect 24254 1187 24255 1232
rect 25598 1187 25599 1232
rect 26846 1187 26847 1232
rect 28190 1187 28191 1232
rect 29438 1187 29439 1232
rect 30686 1187 30687 1232
rect 32030 1187 32031 1232
rect 33278 1187 33279 1232
rect 34526 1187 34527 1232
rect 35294 1187 35295 1232
rect 960 133 961 144
rect 1728 133 1729 144
rect 971 99 972 133
rect 1739 99 1740 133
rect 4382 111 4383 156
rect 5630 111 5631 156
rect 6974 111 6975 156
rect 8222 111 8223 156
rect 9470 111 9471 156
rect 10814 111 10815 156
rect 12062 111 12063 156
rect 12960 133 12961 144
rect 13728 133 13729 144
rect 14496 133 14497 144
rect 12971 99 12972 133
rect 13739 99 13740 133
rect 14507 99 14508 133
rect 15422 111 15423 156
rect 16128 133 16129 144
rect 16139 99 16140 133
rect 17054 111 17055 156
rect 18494 111 18495 156
rect 19488 133 19489 144
rect 20544 133 20545 144
rect 21984 133 21985 144
rect 19499 99 19500 133
rect 20555 99 20556 133
rect 21995 99 21996 133
rect 23006 111 23007 156
rect 24254 111 24255 156
rect 25598 111 25599 156
rect 26846 111 26847 156
rect 28190 111 28191 156
rect 29438 111 29439 156
rect 30686 111 30687 156
rect 32030 111 32031 156
rect 33278 111 33279 156
rect 34526 111 34527 156
<< locali >>
rect 5695 18890 5904 18924
rect 11263 18890 11472 18924
rect 15967 18890 16176 18924
rect 23760 18890 23873 18924
rect 5695 18742 5729 18890
rect 11263 18742 11297 18890
rect 15967 18816 16001 18890
rect 23839 18816 23873 18890
rect 14256 18372 14369 18406
rect 17136 18372 17249 18406
rect 18960 18372 19073 18406
rect 23088 18372 23201 18406
rect 14335 18076 14369 18372
rect 17215 18076 17249 18372
rect 19039 18076 19073 18372
rect 20095 18298 20208 18332
rect 20095 18076 20129 18298
rect 23167 18224 23201 18372
rect 991 17592 1025 17888
rect 2815 17592 2849 17888
rect 5695 17592 5729 17888
rect 7519 17592 7553 17888
rect 991 17558 1104 17592
rect 2815 17558 2928 17592
rect 5695 17558 5808 17592
rect 7519 17558 7632 17592
rect 13663 17000 13697 17222
rect 16543 17000 16577 17222
rect 1488 16966 1601 17000
rect 3312 16966 3425 17000
rect 6192 16966 6305 17000
rect 13584 16966 13697 17000
rect 16464 16966 16577 17000
rect 22416 16966 22625 17000
rect 1567 16818 1601 16966
rect 3391 16818 3425 16966
rect 6271 16744 6305 16966
rect 22591 16818 22625 16966
rect 15967 16334 16001 16482
rect 20095 16334 20129 16556
rect 7519 16300 7632 16334
rect 15967 16300 16080 16334
rect 17791 16300 17904 16334
rect 20095 16300 20208 16334
rect 17791 16078 17825 16300
rect 13471 15634 13584 15668
rect 29599 15634 29712 15668
rect 29599 15412 29633 15634
rect 27295 15002 27329 15076
rect 27216 14968 27329 15002
rect 2640 14894 2753 14928
rect 2719 14746 2753 14894
rect 1951 14410 1985 14558
rect 1951 14376 2064 14410
rect 1951 14228 1985 14376
rect 23952 14228 24065 14262
rect 1471 13596 1505 13892
rect 1951 13596 1985 13892
rect 1471 13562 1584 13596
rect 1872 13562 1985 13596
rect 127 13004 161 13226
rect 31 12970 161 13004
rect 3103 12970 3504 13004
rect 31 12042 65 12970
rect 3103 12748 3137 12970
rect 895 12264 929 12560
rect 1471 12264 1505 12560
rect 2160 12526 2273 12560
rect 29119 12338 29153 12412
rect 29040 12304 29153 12338
rect 895 12230 1008 12264
rect 1471 12230 1584 12264
rect 31 12008 161 12042
rect 127 11786 161 12008
rect 895 11746 929 11820
rect 2047 11746 2081 11894
rect 5695 11746 5729 11894
rect 895 11712 1008 11746
rect 2047 11712 2160 11746
rect 5695 11712 5808 11746
rect 607 10932 641 11228
rect 607 10898 720 10932
rect 1951 10414 1985 10488
rect 720 10380 833 10414
rect 1951 10380 2064 10414
rect 799 10158 833 10380
rect 415 9048 528 9082
rect 816 9048 929 9082
rect 415 8752 449 9048
rect 895 8752 929 9048
rect 816 8234 929 8268
rect 127 7898 161 8120
rect 895 8086 929 8234
rect 1855 8234 1968 8268
rect 1855 8160 1889 8234
rect 31 7864 161 7898
rect 31 5456 65 7864
rect 415 7716 528 7750
rect 415 7420 449 7716
rect 31 5422 161 5456
rect 127 5200 161 5422
rect 31 4978 432 5012
rect 31 2422 65 4978
rect 31 2388 161 2422
rect 127 2166 161 2388
rect 127 1090 161 1460
rect 127 1056 336 1090
rect 19135 350 19169 424
rect 19135 316 19248 350
rect 1392 242 1488 276
rect 14160 242 14256 276
<< metal1 >>
rect 0 20597 36000 20695
rect 7042 20373 12158 20401
rect 7042 20327 7070 20373
rect 4354 20299 4478 20327
rect 4665 20299 4752 20327
rect 6274 20299 6494 20327
rect 6969 20299 7070 20327
rect 34 20225 4286 20253
rect 4258 20179 4286 20225
rect 4834 20225 19646 20253
rect 4834 20179 4862 20225
rect 4258 20151 4862 20179
rect 0 19931 36000 20029
rect 3106 19855 3230 19883
rect 7522 19855 7742 19883
rect 13282 19855 13406 19883
rect 17506 19855 17630 19883
rect 21634 19855 21758 19883
rect 4435 19661 4493 19747
rect 4930 19707 6110 19735
rect 4930 19661 4958 19707
rect 3129 19633 3216 19661
rect 4258 19633 4493 19661
rect 4665 19633 4958 19661
rect 6082 19661 6110 19707
rect 6082 19633 6590 19661
rect 6969 19633 7056 19661
rect 7737 19633 7824 19661
rect 13401 19633 13488 19661
rect 16834 19633 17630 19661
rect 20290 19633 21662 19661
rect 4435 19624 4493 19633
rect 226 19559 2942 19587
rect 226 19439 254 19559
rect 34 19411 254 19439
rect 2914 19439 2942 19559
rect 3394 19559 4094 19587
rect 16834 19559 16862 19633
rect 3394 19439 3422 19559
rect 4066 19513 4094 19559
rect 4066 19485 6014 19513
rect 2914 19411 3422 19439
rect 5986 19439 6014 19485
rect 5986 19411 6206 19439
rect 0 19265 36000 19363
rect 5410 19152 7934 19180
rect 5410 19069 5438 19152
rect 7906 19143 7934 19152
rect 17122 19152 18206 19180
rect 17122 19143 17150 19152
rect 7906 19115 9566 19143
rect 9538 19069 9566 19115
rect 12898 19115 13310 19143
rect 13401 19115 13488 19143
rect 16450 19115 17150 19143
rect 18178 19143 18206 19152
rect 18178 19115 20126 19143
rect 20409 19115 22142 19143
rect 12898 19069 12926 19115
rect 16450 19069 16478 19115
rect 1186 19041 3230 19069
rect 4546 19041 5438 19069
rect 5986 19041 6302 19069
rect 4546 18995 4574 19041
rect 2818 18967 4574 18995
rect 6274 18995 6302 19041
rect 7234 19041 7934 19069
rect 9538 19041 12926 19069
rect 13090 19041 16478 19069
rect 17218 19041 18014 19069
rect 22210 19041 33470 19069
rect 7234 18995 7262 19041
rect 6274 18967 7262 18995
rect 7618 18967 7742 18995
rect 1090 18893 1214 18921
rect 2818 18893 2846 18967
rect 2914 18893 3038 18921
rect 4642 18893 5918 18921
rect 7426 18893 7550 18921
rect 7714 18893 7742 18967
rect 8098 18967 9182 18995
rect 8098 18921 8126 18967
rect 7810 18893 8126 18921
rect 9154 18921 9182 18967
rect 9154 18893 9374 18921
rect 13090 18893 13118 19041
rect 17218 18995 17246 19041
rect 22210 19032 22238 19041
rect 19330 19004 20510 19032
rect 19330 18995 19358 19004
rect 16642 18967 17246 18995
rect 17794 18967 19358 18995
rect 20482 18995 20510 19004
rect 21634 19004 22238 19032
rect 21634 18995 21662 19004
rect 20482 18967 21662 18995
rect 5890 18847 5918 18893
rect 5890 18819 7262 18847
rect 7234 18810 7262 18819
rect 9538 18819 10142 18847
rect 11577 18819 11664 18847
rect 9538 18810 9566 18819
rect 7234 18782 9566 18810
rect 10114 18773 10142 18819
rect 13282 18773 13310 18921
rect 5698 18745 5822 18773
rect 10114 18745 10334 18773
rect 11266 18745 11390 18773
rect 13090 18745 13310 18773
rect 14914 18773 14942 18921
rect 17794 18893 17822 18967
rect 17890 18893 18014 18921
rect 19545 18893 19632 18921
rect 20217 18893 20304 18921
rect 21826 18893 21950 18921
rect 22018 18893 22142 18921
rect 33442 18893 33470 19041
rect 15106 18819 15806 18847
rect 15970 18819 16286 18847
rect 16450 18819 21758 18847
rect 15106 18773 15134 18819
rect 14914 18745 15134 18773
rect 15778 18773 15806 18819
rect 16450 18773 16478 18819
rect 21730 18810 21758 18819
rect 22210 18819 23486 18847
rect 23842 18819 30206 18847
rect 22210 18810 22238 18819
rect 21730 18782 22238 18810
rect 15778 18745 16478 18773
rect 23458 18745 23486 18819
rect 30178 18745 30206 18819
rect 0 18599 36000 18697
rect 34 18523 254 18551
rect 226 18477 254 18523
rect 802 18523 1310 18551
rect 802 18477 830 18523
rect 226 18449 830 18477
rect 1282 18477 1310 18523
rect 7234 18523 7454 18551
rect 21826 18523 22046 18551
rect 7234 18514 7262 18523
rect 1954 18486 7262 18514
rect 22018 18514 22046 18523
rect 26722 18523 26942 18551
rect 22018 18486 26174 18514
rect 1954 18477 1982 18486
rect 26146 18477 26174 18486
rect 26722 18477 26750 18523
rect 1282 18449 1982 18477
rect 15970 18449 16478 18477
rect 26146 18449 26750 18477
rect 15970 18403 15998 18449
rect 2146 18375 3326 18403
rect 3970 18375 4190 18403
rect 4546 18375 6014 18403
rect 5986 18329 6014 18375
rect 6658 18375 6878 18403
rect 8290 18375 8702 18403
rect 12418 18375 15998 18403
rect 16450 18403 16478 18449
rect 16450 18375 19358 18403
rect 21250 18375 22334 18403
rect 6658 18329 6686 18375
rect 1017 18301 1104 18329
rect 2841 18301 2928 18329
rect 4354 18301 4478 18329
rect 4761 18301 4848 18329
rect 5721 18301 5808 18329
rect 5986 18301 6686 18329
rect 7545 18301 7632 18329
rect 9177 18301 9264 18329
rect 9561 18301 9648 18329
rect 11289 18301 11376 18329
rect 13090 18301 13214 18329
rect 16185 18301 16272 18329
rect 17794 18301 17918 18329
rect 1474 18227 1982 18255
rect 1474 18181 1502 18227
rect 1186 18153 1502 18181
rect 1954 18181 1982 18227
rect 1954 18153 3038 18181
rect 5986 18153 7742 18181
rect 11577 18153 13502 18181
rect 14530 18153 15326 18181
rect 16354 18153 18014 18181
rect 14530 18107 14558 18153
rect 14338 18079 14558 18107
rect 15298 18107 15326 18153
rect 15298 18079 15518 18107
rect 17145 18079 17232 18107
rect 18969 18079 19056 18107
rect 19330 18079 19358 18375
rect 21922 18301 22046 18329
rect 22306 18255 22334 18375
rect 22978 18375 25982 18403
rect 22978 18255 23006 18375
rect 25954 18301 25982 18375
rect 22306 18227 23006 18255
rect 23170 18227 29342 18255
rect 20482 18153 22142 18181
rect 20098 18079 20318 18107
rect 0 17933 36000 18031
rect 994 17857 1118 17885
rect 2818 17857 2942 17885
rect 5698 17857 5822 17885
rect 7522 17857 7646 17885
rect 17602 17811 17630 17885
rect 11458 17783 13310 17811
rect 16162 17783 16670 17811
rect 16642 17737 16670 17783
rect 17410 17783 18014 17811
rect 20290 17783 20798 17811
rect 17410 17737 17438 17783
rect 1186 17709 3038 17737
rect 5890 17709 7742 17737
rect 16642 17709 17438 17737
rect 20770 17737 20798 17783
rect 21730 17783 22334 17811
rect 21730 17737 21758 17783
rect 20770 17709 21758 17737
rect 3778 17635 4094 17663
rect 4258 17635 4478 17663
rect 9177 17635 9264 17663
rect 9561 17635 9648 17663
rect 34 17561 3134 17589
rect 3106 17552 3134 17561
rect 4642 17561 5726 17589
rect 11289 17561 11376 17589
rect 12034 17561 12926 17589
rect 13090 17561 13214 17589
rect 13570 17561 14174 17589
rect 16066 17561 16286 17589
rect 17794 17561 17918 17589
rect 18082 17561 18686 17589
rect 4642 17552 4670 17561
rect 3106 17524 4670 17552
rect 5698 17552 5726 17561
rect 5698 17524 6398 17552
rect 6370 17515 6398 17524
rect 6370 17487 7934 17515
rect 7906 17441 7934 17487
rect 12034 17441 12062 17561
rect 12898 17478 12926 17561
rect 13570 17478 13598 17561
rect 14146 17515 14174 17561
rect 18082 17515 18110 17561
rect 14146 17487 14366 17515
rect 12898 17450 13598 17478
rect 1570 17413 2366 17441
rect 3394 17413 4478 17441
rect 6178 17413 6302 17441
rect 7906 17413 8126 17441
rect 11842 17413 12062 17441
rect 13666 17413 13886 17441
rect 14338 17413 14366 17487
rect 16738 17487 18110 17515
rect 18658 17515 18686 17561
rect 19042 17561 19742 17589
rect 20194 17561 20414 17589
rect 21922 17561 22046 17589
rect 22690 17561 24830 17589
rect 18658 17487 18878 17515
rect 16738 17441 16766 17487
rect 19042 17441 19070 17561
rect 16546 17413 16766 17441
rect 18370 17413 19070 17441
rect 19714 17441 19742 17561
rect 20866 17487 21566 17515
rect 20866 17441 20894 17487
rect 19714 17413 19934 17441
rect 20674 17413 20894 17441
rect 21538 17441 21566 17487
rect 22690 17441 22718 17561
rect 21538 17413 21758 17441
rect 22498 17413 22718 17441
rect 24802 17441 24830 17561
rect 24994 17561 28094 17589
rect 24994 17441 25022 17561
rect 28066 17515 28094 17561
rect 28066 17487 28286 17515
rect 24802 17413 25022 17441
rect 28258 17413 28286 17487
rect 0 17267 36000 17365
rect 1282 17191 1694 17219
rect 1666 17071 1694 17191
rect 2818 17191 3326 17219
rect 4834 17191 4958 17219
rect 5986 17191 6398 17219
rect 2818 17071 2846 17191
rect 1666 17043 2846 17071
rect 1209 16969 1296 16997
rect 3033 16969 3120 16997
rect 3874 16923 3902 16997
rect 4089 16969 4176 16997
rect 4258 16969 4862 16997
rect 4930 16969 4958 17191
rect 6370 17145 6398 17191
rect 7426 17191 8030 17219
rect 11650 17191 11966 17219
rect 13090 17191 13694 17219
rect 16258 17191 16574 17219
rect 20505 17191 20592 17219
rect 22306 17191 22430 17219
rect 7426 17145 7454 17191
rect 11938 17182 11966 17191
rect 11938 17154 12638 17182
rect 6370 17117 7454 17145
rect 12610 17145 12638 17154
rect 12610 17117 13598 17145
rect 16377 17117 18302 17145
rect 20290 17117 20798 17145
rect 5218 17043 5726 17071
rect 7618 17043 8030 17071
rect 9250 17043 9374 17071
rect 5218 16997 5246 17043
rect 5026 16969 5246 16997
rect 5698 16997 5726 17043
rect 5698 16969 5918 16997
rect 6850 16969 7742 16997
rect 8002 16969 8030 17043
rect 8217 16969 8304 16997
rect 8386 16969 9182 16997
rect 9346 16969 9374 17043
rect 11458 17043 11966 17071
rect 9634 16969 10334 16997
rect 10425 16969 10512 16997
rect 10594 16969 10910 16997
rect 11458 16969 11486 17043
rect 11554 16969 11774 16997
rect 4258 16923 4286 16969
rect 3778 16895 3902 16923
rect 3970 16895 4286 16923
rect 4834 16849 4862 16969
rect 6082 16895 6686 16923
rect 6082 16849 6110 16895
rect 1186 16821 1598 16849
rect 3010 16821 3422 16849
rect 4834 16821 6110 16849
rect 6658 16849 6686 16895
rect 8386 16849 8414 16969
rect 9154 16923 9182 16969
rect 9634 16923 9662 16969
rect 9154 16895 9662 16923
rect 10306 16923 10334 16969
rect 10594 16923 10622 16969
rect 10306 16895 10622 16923
rect 11938 16923 11966 17043
rect 13186 17043 15806 17071
rect 13186 16923 13214 17043
rect 11938 16895 13214 16923
rect 6658 16821 8414 16849
rect 13378 16849 13406 16997
rect 15778 16969 15806 17043
rect 16834 17043 17054 17071
rect 17890 17043 18110 17071
rect 16834 16997 16862 17043
rect 18082 16997 18110 17043
rect 18466 17043 19742 17071
rect 16258 16969 16862 16997
rect 17986 16923 18014 16997
rect 18082 16969 18302 16997
rect 18466 16923 18494 17043
rect 17986 16895 18494 16923
rect 19714 16923 19742 17043
rect 20290 16969 20318 17117
rect 20770 17071 20798 17117
rect 21730 17117 24350 17145
rect 21730 17071 21758 17117
rect 20770 17043 21758 17071
rect 20386 16969 20606 16997
rect 22210 16969 22814 16997
rect 22786 16923 22814 16969
rect 24418 16969 27710 16997
rect 24418 16923 24446 16969
rect 19714 16895 19934 16923
rect 21922 16895 22238 16923
rect 22786 16895 24446 16923
rect 22210 16849 22238 16895
rect 13378 16821 17918 16849
rect 17890 16812 17918 16821
rect 18562 16821 20990 16849
rect 22210 16821 22622 16849
rect 18562 16812 18590 16821
rect 17890 16784 18590 16812
rect 5890 16747 6302 16775
rect 20962 16747 20990 16821
rect 0 16601 36000 16699
rect 1090 16525 1214 16553
rect 2914 16525 3038 16553
rect 5794 16525 5918 16553
rect 7618 16525 7742 16553
rect 8290 16525 8510 16553
rect 8482 16479 8510 16525
rect 9154 16525 9566 16553
rect 9154 16479 9182 16525
rect 994 16303 1118 16331
rect 3202 16303 3518 16331
rect 3778 16303 3806 16479
rect 8482 16451 9182 16479
rect 3993 16303 4080 16331
rect 6009 16303 6096 16331
rect 6777 16303 6864 16331
rect 6969 16303 7550 16331
rect 3490 16257 3518 16303
rect 3490 16229 3710 16257
rect 8386 16183 8414 16331
rect 8866 16303 9278 16331
rect 9346 16303 9374 16525
rect 9538 16479 9566 16525
rect 10306 16525 10526 16553
rect 11362 16525 11486 16553
rect 13090 16525 13310 16553
rect 16162 16525 16286 16553
rect 17794 16525 18014 16553
rect 19522 16525 20126 16553
rect 20217 16525 20304 16553
rect 21922 16525 22142 16553
rect 10306 16479 10334 16525
rect 9538 16451 10334 16479
rect 11650 16451 12446 16479
rect 12418 16405 12446 16451
rect 13282 16451 13886 16479
rect 13282 16405 13310 16451
rect 12418 16377 13310 16405
rect 13858 16405 13886 16451
rect 15778 16451 15998 16479
rect 24034 16451 24638 16479
rect 15778 16405 15806 16451
rect 24034 16405 24062 16451
rect 13858 16377 15806 16405
rect 17026 16377 24062 16405
rect 24610 16405 24638 16451
rect 24610 16377 30974 16405
rect 9442 16303 9854 16331
rect 9250 16257 9278 16303
rect 9442 16257 9470 16303
rect 9250 16229 9470 16257
rect 9826 16257 9854 16303
rect 10402 16303 11582 16331
rect 10402 16257 10430 16303
rect 9826 16229 10430 16257
rect 11554 16257 11582 16303
rect 12034 16303 12254 16331
rect 13474 16303 13694 16331
rect 22233 16303 22320 16331
rect 24130 16303 24254 16331
rect 24322 16303 24542 16331
rect 30946 16303 30974 16377
rect 12034 16257 12062 16303
rect 11554 16229 12062 16257
rect 6850 16155 8606 16183
rect 18082 16155 22142 16183
rect 22498 16155 23870 16183
rect 22498 16109 22526 16155
rect 17721 16081 17808 16109
rect 21922 16081 22526 16109
rect 23842 16109 23870 16155
rect 23842 16081 24062 16109
rect 0 15935 36000 16033
rect 34 15859 254 15887
rect 226 15739 254 15859
rect 1282 15859 1502 15887
rect 1282 15813 1310 15859
rect 9250 15813 9278 15887
rect 24322 15859 24542 15887
rect 802 15785 1310 15813
rect 3993 15785 4080 15813
rect 8098 15785 8510 15813
rect 8578 15785 9566 15813
rect 10882 15785 11774 15813
rect 24322 15785 24350 15859
rect 802 15739 830 15785
rect 9538 15739 9566 15785
rect 226 15711 830 15739
rect 4930 15711 5342 15739
rect 4930 15665 4958 15711
rect 994 15591 1022 15665
rect 1186 15637 1694 15665
rect 1858 15591 1886 15665
rect 2050 15637 2174 15665
rect 2242 15637 2366 15665
rect 3417 15637 3504 15665
rect 3682 15637 4958 15665
rect 5122 15637 5246 15665
rect 5314 15637 5342 15711
rect 9538 15711 10622 15739
rect 5410 15637 6014 15665
rect 2242 15591 2270 15637
rect 5218 15591 5246 15637
rect 5410 15591 5438 15637
rect 994 15563 1214 15591
rect 994 15489 1022 15563
rect 1186 15517 1214 15563
rect 1666 15563 3614 15591
rect 5218 15563 5438 15591
rect 6178 15591 6206 15665
rect 6681 15637 6768 15665
rect 7042 15591 7070 15665
rect 8217 15637 8304 15665
rect 8482 15637 9470 15665
rect 9538 15637 9566 15711
rect 9634 15637 10046 15665
rect 10594 15637 10622 15711
rect 11746 15665 11774 15785
rect 14722 15711 17918 15739
rect 14722 15665 14750 15711
rect 10690 15637 11678 15665
rect 11746 15637 11870 15665
rect 12153 15637 12240 15665
rect 13401 15637 13488 15665
rect 13666 15637 14750 15665
rect 17890 15665 17918 15711
rect 17890 15637 18110 15665
rect 18201 15637 18288 15665
rect 6178 15563 8222 15591
rect 1666 15517 1694 15563
rect 6178 15517 6206 15563
rect 1186 15489 1694 15517
rect 4546 15489 6206 15517
rect 8194 15517 8222 15563
rect 8482 15517 8510 15637
rect 9442 15591 9470 15637
rect 9634 15591 9662 15637
rect 9442 15563 9662 15591
rect 10018 15591 10046 15637
rect 10690 15591 10718 15637
rect 10018 15563 10718 15591
rect 12418 15563 13214 15591
rect 17913 15563 18000 15591
rect 12418 15517 12446 15563
rect 8194 15489 8510 15517
rect 10882 15489 12446 15517
rect 13186 15517 13214 15563
rect 18754 15517 18782 15665
rect 21849 15637 21936 15665
rect 22306 15637 23006 15665
rect 24034 15637 24350 15665
rect 19138 15563 21662 15591
rect 22137 15563 22224 15591
rect 19138 15517 19166 15563
rect 13186 15489 18782 15517
rect 18946 15489 19166 15517
rect 21634 15517 21662 15563
rect 22306 15517 22334 15637
rect 24898 15591 24926 15665
rect 25113 15637 25200 15665
rect 28848 15637 29054 15665
rect 24898 15563 25022 15591
rect 27106 15563 27600 15591
rect 21634 15489 22334 15517
rect 10882 15480 10910 15489
rect 9250 15452 10910 15480
rect 28258 15452 29438 15480
rect 9250 15443 9278 15452
rect 28258 15443 28286 15452
rect 9058 15415 9278 15443
rect 28066 15415 28286 15443
rect 29410 15443 29438 15452
rect 29410 15415 29630 15443
rect 29721 15415 29808 15443
rect 0 15269 36000 15367
rect 3298 15193 3518 15221
rect 3490 15184 3518 15193
rect 7810 15193 8318 15221
rect 3490 15156 4862 15184
rect 4834 15147 4862 15156
rect 898 15119 2078 15147
rect 4834 15119 6590 15147
rect 898 14999 926 15119
rect 610 14971 926 14999
rect 994 14971 1214 14999
rect 1296 14971 1383 14999
rect 1474 14971 1982 14999
rect 2050 14971 2078 15119
rect 6562 15073 6590 15119
rect 7810 15073 7838 15193
rect 8290 15147 8318 15193
rect 9442 15193 9662 15221
rect 10306 15193 10526 15221
rect 9442 15147 9470 15193
rect 10498 15184 10526 15193
rect 16642 15193 16862 15221
rect 24130 15193 24350 15221
rect 10498 15156 11102 15184
rect 8290 15119 9470 15147
rect 11074 15147 11102 15156
rect 11074 15119 15134 15147
rect 15106 15073 15134 15119
rect 16642 15073 16670 15193
rect 27202 15156 28862 15184
rect 27202 15147 27230 15156
rect 24706 15119 27230 15147
rect 28834 15147 28862 15156
rect 28834 15119 29054 15147
rect 3609 15045 3696 15073
rect 4354 15045 4670 15073
rect 6562 15045 7838 15073
rect 8025 15045 8112 15073
rect 10306 15045 10910 15073
rect 15106 15045 16670 15073
rect 22137 15045 22224 15073
rect 22882 15045 26174 15073
rect 27298 15045 27600 15073
rect 2242 14971 2462 14999
rect 3417 14971 3504 14999
rect 1186 14925 1214 14971
rect 1474 14925 1502 14971
rect 1186 14897 1502 14925
rect 2146 14897 2366 14925
rect 2722 14897 3230 14925
rect 2722 14851 2750 14897
rect 2530 14823 2750 14851
rect 3202 14851 3230 14897
rect 4354 14851 4382 15045
rect 4642 14999 4670 15045
rect 4473 14971 4560 14999
rect 4642 14971 5246 14999
rect 5410 14851 5438 14999
rect 5913 14971 6000 14999
rect 6274 14971 6398 14999
rect 8217 14971 8304 14999
rect 8889 14971 10430 14999
rect 10498 14971 10526 15045
rect 10594 14971 10814 14999
rect 10402 14925 10430 14971
rect 10594 14925 10622 14971
rect 10402 14897 10622 14925
rect 10882 14925 10910 15045
rect 29026 14999 29054 15119
rect 11746 14971 11966 14999
rect 12226 14971 13118 14999
rect 13593 14971 13680 14999
rect 14457 14971 14942 14999
rect 11746 14925 11774 14971
rect 10882 14897 11774 14925
rect 17890 14925 17918 14999
rect 18658 14971 19166 14999
rect 21849 14971 21936 14999
rect 22905 14971 22992 14999
rect 24034 14971 24638 14999
rect 17890 14897 18302 14925
rect 23266 14897 23390 14925
rect 24610 14851 24638 14971
rect 24802 14925 24830 14999
rect 25113 14971 25200 14999
rect 25497 14971 25584 14999
rect 29026 14971 29822 14999
rect 28834 14925 28862 14966
rect 24802 14897 24926 14925
rect 25282 14897 26654 14925
rect 26818 14897 27422 14925
rect 28834 14897 29054 14925
rect 25282 14851 25310 14897
rect 3202 14823 4382 14851
rect 4546 14823 5438 14851
rect 17986 14823 18398 14851
rect 24610 14823 25310 14851
rect 27010 14823 27134 14851
rect 1858 14749 2750 14777
rect 23746 14749 24062 14777
rect 26914 14749 27230 14777
rect 29817 14749 29904 14777
rect 0 14603 36000 14701
rect 514 14527 638 14555
rect 1954 14527 2174 14555
rect 2338 14527 2558 14555
rect 1282 14453 1790 14481
rect 34 14379 350 14407
rect 610 14379 1118 14407
rect 1378 14333 1406 14453
rect 2530 14407 2558 14527
rect 3874 14527 4094 14555
rect 24898 14527 25886 14555
rect 3874 14481 3902 14527
rect 25858 14481 25886 14527
rect 27010 14527 27230 14555
rect 27010 14518 27038 14527
rect 26434 14490 27038 14518
rect 26434 14481 26462 14490
rect 3202 14453 3902 14481
rect 9922 14453 10526 14481
rect 25858 14453 26462 14481
rect 3202 14407 3230 14453
rect 1474 14379 1598 14407
rect 1785 14379 1872 14407
rect 2242 14379 2366 14407
rect 2530 14379 3230 14407
rect 5986 14379 6782 14407
rect 418 14305 542 14333
rect 921 14305 1008 14333
rect 1186 14305 1406 14333
rect 1593 14305 2174 14333
rect 3417 14305 3504 14333
rect 3874 14305 4478 14333
rect 4546 14305 4958 14333
rect 5049 14305 5136 14333
rect 6082 14305 6110 14379
rect 6754 14333 6782 14379
rect 9922 14333 9950 14453
rect 10498 14407 10526 14453
rect 10498 14379 11774 14407
rect 26722 14379 27038 14407
rect 10690 14333 10718 14379
rect 11746 14333 11774 14379
rect 6201 14305 6288 14333
rect 6754 14305 6878 14333
rect 7065 14305 7152 14333
rect 7234 14305 8318 14333
rect 8889 14305 9950 14333
rect 10018 14305 10526 14333
rect 10690 14305 10910 14333
rect 34 14231 254 14259
rect 226 14222 254 14231
rect 1762 14231 1982 14259
rect 3609 14231 3696 14259
rect 226 14194 1214 14222
rect 1186 14185 1214 14194
rect 1762 14185 1790 14231
rect 1186 14157 1790 14185
rect 4450 14185 4478 14305
rect 5218 14231 6014 14259
rect 5218 14185 5246 14231
rect 4450 14157 5246 14185
rect 5986 14185 6014 14231
rect 7234 14185 7262 14305
rect 11554 14259 11582 14333
rect 11746 14305 11966 14333
rect 13593 14305 13680 14333
rect 14553 14305 14640 14333
rect 18201 14305 18288 14333
rect 18946 14305 19166 14333
rect 21849 14305 21936 14333
rect 22905 14305 22992 14333
rect 23266 14305 23774 14333
rect 24610 14305 24926 14333
rect 26626 14305 26942 14333
rect 27010 14305 27038 14379
rect 28848 14305 29054 14333
rect 29817 14305 29904 14333
rect 8025 14231 8112 14259
rect 10978 14231 11870 14259
rect 17913 14231 18000 14259
rect 5986 14157 7262 14185
rect 23746 14185 23774 14305
rect 24034 14231 24254 14259
rect 27394 14231 27600 14259
rect 23746 14157 27038 14185
rect 610 14083 1022 14111
rect 2338 14083 2462 14111
rect 22306 14083 22430 14111
rect 23842 14083 25790 14111
rect 29698 14083 29822 14111
rect 0 13937 36000 14035
rect 1401 13861 1488 13889
rect 1954 13861 2270 13889
rect 26434 13861 26654 13889
rect 10306 13787 10910 13815
rect 10306 13741 10334 13787
rect 3513 13713 3600 13741
rect 8025 13713 8112 13741
rect 8770 13713 10334 13741
rect 10882 13741 10910 13787
rect 11554 13787 12254 13815
rect 11554 13741 11582 13787
rect 10882 13713 11582 13741
rect 8770 13667 8798 13713
rect 12226 13667 12254 13787
rect 24034 13787 24350 13815
rect 24034 13741 24062 13787
rect 24322 13741 24350 13787
rect 17913 13713 18000 13741
rect 23458 13713 24062 13741
rect 24130 13713 24254 13741
rect 24322 13713 24432 13741
rect 27202 13713 27600 13741
rect 441 13639 528 13667
rect 921 13639 1008 13667
rect 1186 13639 1502 13667
rect 1593 13639 1680 13667
rect 2050 13639 2750 13667
rect 2818 13639 2942 13667
rect 3417 13639 3504 13667
rect 3586 13639 4670 13667
rect 5232 13639 5319 13667
rect 2818 13593 2846 13639
rect 3586 13593 3614 13639
rect 130 13565 446 13593
rect 706 13565 1118 13593
rect 2338 13565 2462 13593
rect 2530 13565 3614 13593
rect 4642 13593 4670 13639
rect 5410 13593 5438 13667
rect 4642 13565 5438 13593
rect 610 13417 1310 13445
rect 1689 13417 1776 13445
rect 5986 13417 6014 13667
rect 6105 13639 6782 13667
rect 6864 13639 6951 13667
rect 6754 13593 6782 13639
rect 7138 13593 7166 13667
rect 8217 13639 8798 13667
rect 8889 13639 8990 13667
rect 10425 13639 10512 13667
rect 8962 13593 8990 13639
rect 10786 13593 10814 13667
rect 11673 13639 11760 13667
rect 12057 13639 12144 13667
rect 12226 13639 13694 13667
rect 14553 13639 14640 13667
rect 18201 13639 18288 13667
rect 6754 13565 8414 13593
rect 8962 13565 10814 13593
rect 18946 13593 18974 13667
rect 21849 13639 21936 13667
rect 22905 13639 22992 13667
rect 23961 13639 24048 13667
rect 24610 13639 24926 13667
rect 28848 13639 29054 13667
rect 29698 13639 29904 13667
rect 18946 13565 19070 13593
rect 23577 13565 23664 13593
rect 23746 13565 23870 13593
rect 8386 13519 8414 13565
rect 8386 13491 8894 13519
rect 22306 13491 22430 13519
rect 8866 13482 8894 13491
rect 8866 13454 9662 13482
rect 9634 13445 9662 13454
rect 9634 13417 9854 13445
rect 23842 13417 24158 13445
rect 0 13271 36000 13369
rect 34 13195 158 13223
rect 17986 13149 18014 13223
rect 21730 13195 21950 13223
rect 21922 13186 21950 13195
rect 24802 13195 25022 13223
rect 21922 13158 22622 13186
rect 22594 13149 22622 13158
rect 24802 13149 24830 13195
rect 17986 13121 18398 13149
rect 22594 13121 24830 13149
rect 322 13047 446 13075
rect 706 13047 830 13075
rect 1186 13047 2078 13075
rect 1186 13001 1214 13047
rect 441 12973 528 13001
rect 898 12927 926 13001
rect 1090 12973 1214 13001
rect 1378 12927 1406 13001
rect 1570 12973 1598 13047
rect 2050 13001 2078 13047
rect 2242 13047 3230 13075
rect 2242 13001 2270 13047
rect 1858 12927 1886 13001
rect 2050 12973 2270 13001
rect 706 12899 926 12927
rect 1282 12899 1886 12927
rect 3202 12927 3230 13047
rect 4930 13047 5342 13075
rect 4930 13001 4958 13047
rect 3417 12973 3504 13001
rect 4546 12973 4958 13001
rect 5136 12973 5223 13001
rect 5314 12973 5342 13047
rect 6466 13047 6878 13075
rect 22329 13047 22416 13075
rect 25570 13047 25694 13075
rect 25762 13047 26750 13075
rect 6466 13001 6494 13047
rect 5913 12973 6000 13001
rect 6178 12973 6494 13001
rect 6585 12973 6672 13001
rect 6850 12973 6878 13047
rect 25570 13005 25598 13047
rect 8217 12973 8304 13001
rect 8889 12973 8976 13001
rect 9058 12973 9470 13001
rect 9753 12973 10526 13001
rect 10905 12973 10992 13001
rect 11673 12973 11760 13001
rect 12057 12973 12144 13001
rect 13593 12973 13680 13001
rect 14553 12973 14640 13001
rect 18201 12973 18782 13001
rect 18946 12973 19166 13001
rect 21849 12973 21936 13001
rect 22905 12973 22992 13001
rect 23938 12973 24254 13001
rect 25858 12973 25982 13001
rect 29698 12973 29904 13001
rect 3202 12899 3614 12927
rect 8025 12899 8112 12927
rect 18754 12853 18782 12973
rect 19234 12899 24158 12927
rect 25680 12899 26270 12927
rect 29602 12899 29808 12927
rect 19234 12853 19262 12899
rect 2434 12825 2942 12853
rect 18754 12825 19262 12853
rect 23554 12825 26654 12853
rect 2434 12816 2462 12825
rect 1858 12788 2462 12816
rect 1858 12779 1886 12788
rect 1666 12751 1886 12779
rect 2914 12779 2942 12825
rect 2914 12751 3134 12779
rect 27321 12751 27408 12779
rect 0 12605 36000 12703
rect 34 12529 254 12557
rect 226 12483 254 12529
rect 706 12529 926 12557
rect 1401 12529 1488 12557
rect 706 12483 734 12529
rect 2050 12483 2078 12557
rect 2242 12529 4382 12557
rect 4354 12520 4382 12529
rect 5794 12529 6686 12557
rect 24034 12529 24254 12557
rect 26818 12529 27038 12557
rect 5794 12520 5822 12529
rect 4354 12492 5822 12520
rect 226 12455 734 12483
rect 1570 12455 2654 12483
rect 322 12307 1982 12335
rect 2626 12307 2654 12455
rect 3202 12418 4190 12446
rect 3202 12409 3230 12418
rect 3010 12381 3230 12409
rect 4162 12409 4190 12418
rect 4162 12381 5438 12409
rect 3010 12335 3038 12381
rect 2745 12307 3038 12335
rect 3129 12307 3216 12335
rect 3298 12261 3326 12335
rect 3490 12307 3614 12335
rect 3778 12261 3806 12335
rect 130 12233 446 12261
rect 633 12233 720 12261
rect 1209 12233 1296 12261
rect 1689 12233 1776 12261
rect 1872 12233 1959 12261
rect 2050 12233 2174 12261
rect 3298 12233 3806 12261
rect 4258 12261 4286 12335
rect 4354 12307 4382 12381
rect 4642 12261 4670 12335
rect 4834 12307 4862 12381
rect 5218 12261 5246 12335
rect 5410 12307 5438 12381
rect 5602 12307 6110 12335
rect 6178 12307 6494 12335
rect 6658 12307 6686 12529
rect 22594 12455 27422 12483
rect 7234 12381 7742 12409
rect 7234 12335 7262 12381
rect 4258 12233 5246 12261
rect 6466 12261 6494 12307
rect 6850 12261 6878 12335
rect 7042 12307 7262 12335
rect 7330 12261 7358 12335
rect 7714 12307 7742 12381
rect 10786 12381 11006 12409
rect 7906 12307 8414 12335
rect 8962 12307 9278 12335
rect 9753 12307 10718 12335
rect 10786 12307 10814 12381
rect 7906 12261 7934 12307
rect 6466 12233 7934 12261
rect 10690 12261 10718 12307
rect 11074 12261 11102 12335
rect 11673 12307 11760 12335
rect 12057 12307 12144 12335
rect 14146 12307 14270 12335
rect 14553 12307 14640 12335
rect 22594 12307 22622 12455
rect 24130 12381 24336 12409
rect 29122 12381 29808 12409
rect 23458 12307 23582 12335
rect 25584 12307 25790 12335
rect 25954 12307 28478 12335
rect 29698 12307 29904 12335
rect 10690 12233 11102 12261
rect 14146 12233 14174 12307
rect 24130 12233 26174 12261
rect 28569 12233 28656 12261
rect 28834 12233 29630 12261
rect 3298 12159 3326 12233
rect 537 12085 624 12113
rect 1186 12085 1886 12113
rect 23193 12085 23280 12113
rect 26050 12085 26174 12113
rect 27490 12085 27710 12113
rect 28738 12085 28862 12113
rect 0 11939 36000 12037
rect 1186 11863 1502 11891
rect 1666 11863 1886 11891
rect 1977 11863 2064 11891
rect 2338 11863 4766 11891
rect 4738 11854 4766 11863
rect 5506 11863 5726 11891
rect 23170 11863 23390 11891
rect 24130 11863 25886 11891
rect 5506 11854 5534 11863
rect 4738 11826 5534 11854
rect 130 11789 926 11817
rect 1090 11743 1118 11817
rect 1954 11789 2654 11817
rect 2626 11780 2654 11789
rect 4354 11789 4574 11817
rect 4354 11780 4382 11789
rect 2626 11752 4382 11780
rect 4546 11743 4574 11789
rect 6178 11743 6206 11817
rect 25570 11789 26942 11817
rect 27106 11743 27134 11891
rect 34 11715 446 11743
rect 633 11715 720 11743
rect 1090 11715 1310 11743
rect 1497 11715 1584 11743
rect 2338 11715 2462 11743
rect 4546 11715 5150 11743
rect 5986 11715 8030 11743
rect 514 11641 2270 11669
rect 2338 11641 2750 11669
rect 2841 11641 2928 11669
rect 3225 11641 3312 11669
rect 3417 11641 3504 11669
rect 4258 11641 4382 11669
rect 4546 11641 4766 11669
rect 5122 11641 5150 11715
rect 5241 11641 5328 11669
rect 6082 11641 6206 11669
rect 6370 11641 6398 11715
rect 6969 11641 7070 11669
rect 7234 11641 7262 11715
rect 2338 11558 2366 11641
rect 7042 11595 7070 11641
rect 7810 11595 7838 11669
rect 8002 11641 8030 11715
rect 8962 11715 9182 11743
rect 8962 11669 8990 11715
rect 9154 11669 9182 11715
rect 10210 11715 14462 11743
rect 22786 11715 22910 11743
rect 23266 11715 23486 11743
rect 26338 11715 27134 11743
rect 10210 11669 10238 11715
rect 11074 11669 11102 11715
rect 8290 11641 8990 11669
rect 9058 11595 9086 11669
rect 9154 11641 9662 11669
rect 9826 11641 10238 11669
rect 10905 11641 10992 11669
rect 11074 11641 11198 11669
rect 11673 11641 11774 11669
rect 12130 11641 12158 11715
rect 802 11530 2366 11558
rect 802 11521 830 11530
rect 610 11493 830 11521
rect 2530 11493 5438 11521
rect 2530 11447 2558 11493
rect 706 11419 2558 11447
rect 5410 11447 5438 11493
rect 5602 11447 5630 11595
rect 7042 11567 7838 11595
rect 8866 11567 9086 11595
rect 11746 11595 11774 11641
rect 13186 11595 13214 11669
rect 13570 11641 13598 11715
rect 14434 11669 14462 11715
rect 14338 11595 14366 11669
rect 14434 11641 14942 11669
rect 25584 11641 25790 11669
rect 25954 11641 26174 11669
rect 27417 11641 27504 11669
rect 11746 11567 14366 11595
rect 24034 11567 24336 11595
rect 25762 11493 25790 11641
rect 28642 11595 28670 11743
rect 29698 11641 29904 11669
rect 27010 11567 27230 11595
rect 28642 11567 29808 11595
rect 5410 11419 5630 11447
rect 26050 11419 26174 11447
rect 27490 11419 27710 11447
rect 0 11273 36000 11371
rect 130 11197 638 11225
rect 994 11197 1214 11225
rect 1378 11197 1790 11225
rect 1762 11151 1790 11197
rect 6850 11197 7070 11225
rect 24034 11197 24158 11225
rect 26937 11197 27024 11225
rect 4066 11160 5054 11188
rect 4066 11151 4094 11160
rect 1497 11123 1584 11151
rect 1762 11123 4094 11151
rect 5026 11077 5054 11160
rect 6850 11151 6878 11197
rect 5794 11123 6878 11151
rect 14146 11123 14366 11151
rect 5794 11077 5822 11123
rect 4258 11049 4670 11077
rect 5026 11049 5822 11077
rect 802 10975 2270 11003
rect 34 10855 62 10929
rect 921 10901 1008 10929
rect 1090 10855 1118 10929
rect 1282 10901 1406 10929
rect 2073 10901 2160 10929
rect 2338 10901 2462 10929
rect 34 10827 1118 10855
rect 3202 10855 3230 11003
rect 3298 10975 3518 11003
rect 3609 10975 3696 11003
rect 3490 10929 3518 10975
rect 3778 10929 3806 11003
rect 4258 10975 4286 11049
rect 4354 10929 4382 11003
rect 4642 10975 4670 11049
rect 4834 10929 4862 11003
rect 6009 10975 6096 11003
rect 6274 10975 6398 11003
rect 7042 10975 7166 11003
rect 7714 10975 9086 11003
rect 9154 10975 10238 11003
rect 10786 10975 11966 11003
rect 12249 10975 12336 11003
rect 13017 10975 13104 11003
rect 13666 10975 14270 11003
rect 14338 10975 14366 11123
rect 23650 11049 24336 11077
rect 28834 11049 29808 11077
rect 14434 10975 14654 11003
rect 25584 10975 25790 11003
rect 26073 10975 26160 11003
rect 26242 10975 26366 11003
rect 27417 10975 27504 11003
rect 29698 10975 29904 11003
rect 3490 10901 4862 10929
rect 14242 10929 14270 10975
rect 14434 10929 14462 10975
rect 14242 10901 14462 10929
rect 23458 10901 23678 10929
rect 3202 10827 3326 10855
rect 2338 10753 3134 10781
rect 26073 10753 26160 10781
rect 27490 10753 27614 10781
rect 0 10607 36000 10705
rect 34 10457 2174 10485
rect 13090 10457 13790 10485
rect 13090 10411 13118 10457
rect 226 10383 446 10411
rect 2050 10383 2846 10411
rect 3010 10383 3134 10411
rect 3202 10383 8414 10411
rect 514 10309 1022 10337
rect 1113 10309 1200 10337
rect 1378 10309 2174 10337
rect 3298 10309 3422 10337
rect 3586 10309 3614 10383
rect 4258 10309 4382 10337
rect 4450 10309 4478 10383
rect 5145 10309 5232 10337
rect 5314 10309 5342 10383
rect 5986 10309 6110 10337
rect 6466 10309 6494 10383
rect 8386 10337 8414 10383
rect 9826 10383 13118 10411
rect 9826 10337 9854 10383
rect 10018 10337 10046 10383
rect 11458 10337 11486 10383
rect 12898 10337 12926 10383
rect 13762 10337 13790 10457
rect 26146 10341 26174 10485
rect 8217 10309 8304 10337
rect 8386 10309 9854 10337
rect 994 10263 1022 10309
rect 4258 10263 4286 10309
rect 994 10235 1118 10263
rect 2338 10235 3230 10263
rect 3202 10189 3230 10235
rect 3682 10235 4286 10263
rect 9922 10263 9950 10337
rect 10018 10309 10238 10337
rect 11266 10263 11294 10337
rect 11458 10309 11678 10337
rect 12802 10263 12830 10337
rect 12898 10309 13118 10337
rect 13570 10263 13598 10337
rect 13762 10309 14078 10337
rect 25584 10309 25790 10337
rect 27490 10309 27696 10337
rect 25762 10263 25790 10309
rect 9922 10235 11390 10263
rect 12802 10235 13598 10263
rect 17890 10235 21950 10263
rect 23842 10235 24336 10263
rect 25762 10235 25968 10263
rect 28944 10235 29054 10263
rect 3682 10189 3710 10235
rect 802 10161 926 10189
rect 1282 10161 1790 10189
rect 3202 10161 3710 10189
rect 1282 10115 1310 10161
rect 706 10087 1310 10115
rect 1762 10115 1790 10161
rect 1762 10087 1982 10115
rect 0 9941 36000 10039
rect 17218 9865 17438 9893
rect 802 9791 3326 9819
rect 8578 9791 9278 9819
rect 8578 9745 8606 9791
rect 3394 9717 3902 9745
rect 3394 9671 3422 9717
rect 3874 9671 3902 9717
rect 8002 9717 8606 9745
rect 9250 9745 9278 9791
rect 11170 9791 11774 9819
rect 11170 9745 11198 9791
rect 9250 9717 11198 9745
rect 11746 9745 11774 9791
rect 17410 9745 17438 9865
rect 19522 9865 19742 9893
rect 19522 9745 19550 9865
rect 11746 9717 13022 9745
rect 17410 9717 19550 9745
rect 8002 9671 8030 9717
rect 537 9643 1502 9671
rect 1954 9643 2174 9671
rect 2146 9597 2174 9643
rect 2914 9643 3134 9671
rect 3298 9643 3422 9671
rect 2914 9597 2942 9643
rect 3586 9597 3614 9671
rect 34 9569 542 9597
rect 802 9569 1118 9597
rect 2146 9569 2942 9597
rect 3490 9569 3614 9597
rect 3682 9643 3806 9671
rect 3874 9643 4286 9671
rect 4834 9643 6014 9671
rect 6393 9643 6480 9671
rect 7618 9643 8030 9671
rect 8112 9643 8199 9671
rect 34 9495 62 9569
rect 3682 9523 3710 9643
rect 7618 9569 7646 9643
rect 8674 9597 8702 9671
rect 9072 9643 9159 9671
rect 11289 9643 11390 9671
rect 11577 9643 11664 9671
rect 11362 9597 11390 9643
rect 8674 9569 11390 9597
rect 8674 9523 8702 9569
rect 3298 9495 3710 9523
rect 7906 9495 8702 9523
rect 0 9275 36000 9373
rect 706 9199 926 9227
rect 898 9079 926 9199
rect 3010 9199 3710 9227
rect 3010 9079 3038 9199
rect 3970 9125 4670 9153
rect 3970 9079 3998 9125
rect 898 9051 3038 9079
rect 3490 9051 3998 9079
rect 3490 9005 3518 9051
rect 322 8977 638 9005
rect 3202 8931 3230 9005
rect 3298 8977 3518 9005
rect 3586 8931 3614 9005
rect 3778 8977 3806 9051
rect 4642 9005 4670 9125
rect 5698 9125 6302 9153
rect 5698 9005 5726 9125
rect 6274 9079 6302 9125
rect 7906 9125 8990 9153
rect 6274 9051 7070 9079
rect 7042 9005 7070 9051
rect 7906 9005 7934 9125
rect 8962 9005 8990 9125
rect 4258 8977 4478 9005
rect 4642 8977 5726 9005
rect 5986 8977 6686 9005
rect 7042 8977 7934 9005
rect 8217 8977 8798 9005
rect 8962 8977 10046 9005
rect 10233 8977 10320 9005
rect 3202 8903 3614 8931
rect 1282 8783 1310 8857
rect 4450 8829 7742 8857
rect 4450 8783 4478 8829
rect 130 8755 446 8783
rect 898 8755 1310 8783
rect 4258 8755 4478 8783
rect 7714 8783 7742 8829
rect 7714 8755 7934 8783
rect 0 8609 36000 8707
rect 802 8533 1022 8561
rect 994 8487 1022 8533
rect 1570 8533 2078 8561
rect 2530 8533 2846 8561
rect 1570 8487 1598 8533
rect 994 8459 1598 8487
rect 2530 8413 2558 8533
rect 6274 8459 6974 8487
rect 1762 8385 2558 8413
rect 2626 8385 3614 8413
rect 418 8311 2462 8339
rect 2530 8265 2558 8385
rect 226 8237 542 8265
rect 1378 8237 2270 8265
rect 2338 8191 2366 8265
rect 2530 8237 2654 8265
rect 34 8163 2366 8191
rect 3202 8191 3230 8339
rect 3298 8311 3518 8339
rect 3586 8311 3614 8385
rect 6274 8339 6302 8459
rect 6946 8413 6974 8459
rect 7426 8459 8126 8487
rect 7426 8413 7454 8459
rect 6946 8385 7454 8413
rect 8098 8413 8126 8459
rect 8098 8385 8894 8413
rect 3490 8265 3518 8311
rect 3778 8265 3806 8339
rect 5913 8311 6302 8339
rect 6393 8311 6878 8339
rect 7545 8311 7632 8339
rect 7810 8311 8030 8339
rect 8866 8311 8894 8385
rect 9058 8311 9278 8339
rect 3490 8237 3806 8265
rect 6850 8265 6878 8311
rect 7810 8265 7838 8311
rect 9058 8265 9086 8311
rect 6850 8237 9086 8265
rect 3202 8163 3518 8191
rect 130 8089 926 8117
rect 2146 8089 2270 8117
rect 0 7943 36000 8041
rect 7618 7793 8894 7821
rect 802 7719 1022 7747
rect 2242 7719 3038 7747
rect 3202 7719 3422 7747
rect 322 7645 638 7673
rect 3394 7645 3422 7719
rect 7810 7719 7934 7747
rect 3490 7599 3518 7673
rect 5410 7645 5918 7673
rect 6274 7645 7742 7673
rect 7810 7645 7838 7719
rect 7906 7645 8126 7673
rect 8866 7645 8894 7793
rect 9058 7645 9278 7673
rect 802 7571 3518 7599
rect 7714 7599 7742 7645
rect 7906 7599 7934 7645
rect 9058 7599 9086 7645
rect 7714 7571 9182 7599
rect 15778 7571 17630 7599
rect 226 7423 446 7451
rect 0 7277 36000 7375
rect 1570 7201 1790 7229
rect 5314 7127 6110 7155
rect 5314 7081 5342 7127
rect 3490 7053 5342 7081
rect 3490 7007 3518 7053
rect 322 6979 638 7007
rect 1570 6979 1790 7007
rect 3202 6933 3230 7007
rect 3298 6979 3518 7007
rect 3586 6933 3614 7007
rect 3778 6979 3806 7053
rect 6082 7007 6110 7127
rect 5410 6979 5918 7007
rect 6082 6979 6302 7007
rect 7906 6979 8798 7007
rect 9081 6979 9168 7007
rect 130 6905 542 6933
rect 802 6905 1214 6933
rect 3202 6905 3614 6933
rect 706 6757 1598 6785
rect 0 6611 36000 6709
rect 706 6535 1406 6563
rect 2242 6387 3134 6415
rect 2242 6341 2270 6387
rect 322 6313 446 6341
rect 2050 6313 2270 6341
rect 3106 6341 3134 6387
rect 3106 6313 3326 6341
rect 3417 6313 3504 6341
rect 610 6239 1886 6267
rect 610 6193 638 6239
rect 34 6165 638 6193
rect 1858 6193 1886 6239
rect 1858 6165 4286 6193
rect 0 5945 36000 6043
rect 706 5869 1214 5897
rect 1762 5721 2942 5749
rect 1762 5675 1790 5721
rect 130 5647 446 5675
rect 1570 5647 1790 5675
rect 2914 5675 2942 5721
rect 3490 5721 3710 5749
rect 3490 5675 3518 5721
rect 3682 5675 3710 5721
rect 2914 5647 3230 5675
rect 3298 5647 3518 5675
rect 3202 5601 3230 5647
rect 3586 5601 3614 5675
rect 3682 5647 3806 5675
rect 610 5573 1406 5601
rect 3202 5573 3614 5601
rect 3970 5573 5822 5601
rect 610 5527 638 5573
rect 34 5499 638 5527
rect 1378 5527 1406 5573
rect 3970 5527 3998 5573
rect 1378 5499 3134 5527
rect 3106 5490 3134 5499
rect 3778 5499 3998 5527
rect 5794 5527 5822 5573
rect 5794 5499 6014 5527
rect 3778 5490 3806 5499
rect 3106 5462 3806 5490
rect 0 5279 36000 5377
rect 130 5203 542 5231
rect 226 4907 5246 4935
rect 226 4861 254 4907
rect 34 4833 254 4861
rect 5218 4861 5246 4907
rect 5218 4833 5438 4861
rect 0 4613 36000 4711
rect 921 4537 1008 4565
rect 4066 4343 4094 4417
rect 825 4315 912 4343
rect 4066 4315 11774 4343
rect 11746 4241 11774 4315
rect 0 3947 36000 4045
rect 1570 3723 2078 3751
rect 1209 3575 1296 3603
rect 0 3281 36000 3379
rect 1186 2983 1310 3011
rect 514 2909 1886 2937
rect 994 2761 1118 2789
rect 1858 2761 1982 2789
rect 0 2615 36000 2713
rect 1785 2539 1872 2567
rect 1977 2539 2064 2567
rect 34 2465 350 2493
rect 514 2391 1022 2419
rect 3033 2391 3120 2419
rect 1282 2317 1886 2345
rect 16834 2317 16958 2345
rect 2073 2243 2160 2271
rect 15490 2243 22334 2271
rect 34 2169 158 2197
rect 22306 2169 22334 2243
rect 1017 2095 1104 2123
rect 2818 2095 2942 2123
rect 17337 2095 17424 2123
rect 0 1949 36000 2047
rect 1785 1873 1872 1901
rect 16930 1873 18398 1901
rect 514 1651 1118 1679
rect 1881 1651 1968 1679
rect 13858 1605 13886 1679
rect 13968 1651 14055 1679
rect 16066 1651 16190 1679
rect 17026 1651 17438 1679
rect 17794 1651 18302 1679
rect 1282 1577 1886 1605
rect 3298 1577 3902 1605
rect 13858 1577 21758 1605
rect 16258 1503 17630 1531
rect 130 1429 1118 1457
rect 2338 1429 2654 1457
rect 3129 1429 3216 1457
rect 14242 1429 14558 1457
rect 16834 1429 16958 1457
rect 0 1283 36000 1381
rect 1785 1207 1872 1235
rect 2050 1207 2174 1235
rect 3801 1207 3888 1235
rect 13762 1207 13982 1235
rect 15993 1207 16080 1235
rect 18274 1207 18398 1235
rect 19714 1087 19742 1161
rect 1282 1059 2366 1087
rect 2530 1059 3998 1087
rect 13954 1059 14270 1087
rect 14530 1059 15422 1087
rect 16185 1059 16272 1087
rect 16930 1059 17726 1087
rect 19714 1059 32894 1087
rect 2530 1013 2558 1059
rect 130 985 2558 1013
rect 2626 985 3614 1013
rect 13186 985 13406 1013
rect 14722 985 16862 1013
rect 226 911 1598 939
rect 2146 911 2750 939
rect 2818 911 3422 939
rect 3490 911 3806 939
rect 226 865 254 911
rect 34 837 254 865
rect 1570 865 1598 911
rect 20002 865 20030 939
rect 33058 911 33854 939
rect 33058 865 33086 911
rect 1570 837 1790 865
rect 20002 837 33086 865
rect 33826 865 33854 911
rect 33826 837 34046 865
rect 921 763 1008 791
rect 15225 763 15312 791
rect 0 617 36000 715
rect 3394 541 3518 569
rect 9730 541 9950 569
rect 9922 495 9950 541
rect 12418 541 12638 569
rect 13305 541 13392 569
rect 12418 495 12446 541
rect 9922 467 12446 495
rect 19042 467 31838 495
rect 31810 421 31838 467
rect 35746 467 35966 495
rect 35746 421 35774 467
rect 2626 393 2750 421
rect 2818 393 2942 421
rect 3033 393 3120 421
rect 3216 393 3303 421
rect 6274 393 9566 421
rect 14914 393 15710 421
rect 16546 393 19166 421
rect 6274 347 6302 393
rect 802 319 1022 347
rect 1762 319 2174 347
rect 3010 199 3038 347
rect 3778 319 3902 347
rect 6082 319 6302 347
rect 9538 347 9566 393
rect 15682 347 15710 393
rect 25282 347 25310 421
rect 31810 393 35774 421
rect 9538 319 12830 347
rect 13570 319 15326 347
rect 15682 319 15902 347
rect 19906 319 20126 347
rect 20962 319 21566 347
rect 22402 319 25310 347
rect 20098 273 20126 319
rect 21538 273 21566 319
rect 3202 245 5918 273
rect 3202 199 3230 245
rect 3010 171 3230 199
rect 5890 199 5918 245
rect 18850 199 18878 273
rect 20098 245 20318 273
rect 21538 245 21758 273
rect 25474 245 31646 273
rect 25474 199 25502 245
rect 5890 171 14270 199
rect 14338 171 18494 199
rect 18850 171 25502 199
rect 31618 199 31646 245
rect 31618 171 31838 199
rect 0 -49 36000 49
<< metal2 >>
rect 0 20595 97 20623
rect 34 20225 62 20595
rect 0 20077 97 20105
rect 34 19787 62 20077
rect 3106 19855 3134 20646
rect 4450 19707 4478 20646
rect 0 19633 97 19661
rect 34 19411 62 19633
rect 0 19115 97 19143
rect 34 18811 62 19115
rect 1282 18921 1310 19069
rect 3202 19041 3230 19661
rect 4258 19217 4286 19661
rect 4738 19439 4766 20327
rect 5026 19513 5054 19815
rect 6274 19633 6302 20327
rect 7042 19633 7070 20327
rect 7522 19855 7550 20646
rect 5026 19485 5150 19513
rect 4738 19411 4862 19439
rect 4258 19189 4382 19217
rect 0 18671 97 18699
rect 34 18523 62 18671
rect 0 18153 97 18181
rect 34 17835 62 18153
rect 1090 17737 1118 18921
rect 1282 18893 1406 18921
rect 1378 18329 1406 18893
rect 0 17709 97 17737
rect 994 17709 1118 17737
rect 1282 18301 1406 18329
rect 34 17561 62 17709
rect 0 17191 97 17219
rect 34 17103 62 17191
rect 994 16997 1022 17709
rect 1282 17191 1310 18301
rect 994 16969 1118 16997
rect 1090 16849 1118 16969
rect 1090 16821 1214 16849
rect 0 16747 97 16775
rect 34 16493 62 16747
rect 1090 16525 1118 16821
rect 0 16229 97 16257
rect 34 15859 62 16229
rect 0 15785 97 15813
rect 34 15591 62 15785
rect 34 15563 350 15591
rect 0 15267 97 15295
rect 34 14925 62 15267
rect 34 14897 158 14925
rect 0 14823 97 14851
rect 34 14379 62 14823
rect 130 14777 158 14897
rect 130 14749 206 14777
rect 0 14305 97 14333
rect 34 14231 62 14305
rect 0 13861 97 13889
rect 34 13519 62 13861
rect 178 13741 206 14749
rect 130 13713 206 13741
rect 130 13565 158 13713
rect 34 13491 158 13519
rect 0 13417 97 13445
rect 34 13195 62 13417
rect 130 13371 158 13491
rect 130 13343 206 13371
rect 0 12899 97 12927
rect 34 12529 62 12899
rect 0 12455 97 12483
rect 34 12345 62 12455
rect 178 12409 206 13343
rect 322 13047 350 15563
rect 610 14527 638 14999
rect 514 14254 542 14333
rect 994 14305 1022 16331
rect 1282 16127 1310 16997
rect 1474 15665 1502 15887
rect 1186 15591 1214 15665
rect 1474 15637 1598 15665
rect 1186 15563 1310 15591
rect 1282 14453 1310 15563
rect 1570 15147 1598 15637
rect 1474 15119 1598 15147
rect 2050 15119 2078 15665
rect 1090 14379 1214 14407
rect 514 13001 542 13715
rect 994 13639 1022 14111
rect 1090 13445 1118 13593
rect 1042 13417 1118 13445
rect 130 12381 206 12409
rect 322 12973 542 13001
rect 130 12233 158 12381
rect 322 12307 350 12973
rect 802 12779 830 13075
rect 1042 12779 1070 13417
rect 1186 12853 1214 14379
rect 1474 13861 1502 15119
rect 1666 14971 2270 14999
rect 1282 12899 1310 13445
rect 1186 12825 1310 12853
rect 802 12751 926 12779
rect 1042 12751 1118 12779
rect 898 12557 926 12751
rect 706 12529 926 12557
rect 0 11937 97 11965
rect 34 11715 62 11937
rect 0 11493 97 11521
rect 610 11493 638 12113
rect 706 11743 734 12529
rect 706 11715 830 11743
rect 34 11225 62 11493
rect 802 11447 830 11715
rect 898 11641 926 12335
rect 802 11419 926 11447
rect 898 11225 926 11419
rect 34 11197 158 11225
rect 802 11197 926 11225
rect 802 11077 830 11197
rect 1090 11151 1118 12751
rect 706 11049 830 11077
rect 994 11123 1118 11151
rect 0 10975 97 11003
rect 34 10901 62 10975
rect 0 10531 97 10559
rect 34 10457 62 10531
rect 34 10041 62 10177
rect 0 10013 97 10041
rect 226 9819 254 10411
rect 706 10337 734 11049
rect 706 10309 830 10337
rect 802 10189 830 10309
rect 994 10263 1022 11123
rect 1172 11102 1228 11243
rect 1186 10271 1214 10337
rect 994 10235 1070 10263
rect 802 10161 926 10189
rect 34 9791 254 9819
rect 34 9597 62 9791
rect 0 9569 97 9597
rect 34 9079 62 9523
rect 0 9051 97 9079
rect 34 8755 158 8783
rect 34 8635 62 8755
rect 0 8607 97 8635
rect 322 8561 350 9005
rect 610 8977 638 9671
rect 898 8561 926 10161
rect 1042 9745 1070 10235
rect 1042 9717 1118 9745
rect 1090 8931 1118 9717
rect 1282 9523 1310 12825
rect 1474 12529 1502 13667
rect 1666 13639 1694 14971
rect 1858 13519 1886 14777
rect 2146 14527 2174 14925
rect 2338 14527 2366 17441
rect 2914 16849 2942 18921
rect 3298 17071 3326 18403
rect 4162 18323 4190 18403
rect 4354 18107 4382 19189
rect 4546 18375 4574 18839
rect 4258 18079 4382 18107
rect 3298 17043 3422 17071
rect 2914 16821 3038 16849
rect 2914 16525 2942 16821
rect 3106 16331 3134 16997
rect 3010 16303 3134 16331
rect 1858 13491 1934 13519
rect 1570 12409 1598 12483
rect 1474 12381 1598 12409
rect 1474 11863 1502 12381
rect 1666 11863 1694 12779
rect 1762 12233 1790 13445
rect 1906 12779 1934 13491
rect 1906 12751 1982 12779
rect 1954 12483 1982 12751
rect 2050 12529 2078 13667
rect 2242 13149 2270 14407
rect 2434 13565 2462 14111
rect 2242 13121 2366 13149
rect 1954 12455 2078 12483
rect 1858 12261 1886 12373
rect 1858 12233 1982 12261
rect 1858 11817 1886 12113
rect 1954 11965 1982 12233
rect 2050 12039 2078 12455
rect 2338 12187 2366 13121
rect 2242 12159 2366 12187
rect 2050 12011 2174 12039
rect 1954 11937 2078 11965
rect 2050 11863 2078 11937
rect 1858 11789 1982 11817
rect 1474 9643 1502 11669
rect 1570 11123 1598 11743
rect 2146 11669 2174 12011
rect 2242 11965 2270 12159
rect 2818 12113 2846 12335
rect 3010 12187 3038 16303
rect 3394 16257 3422 17043
rect 3778 16451 3806 17663
rect 4258 17071 4286 18079
rect 4450 17413 4478 17497
rect 4834 17191 4862 19411
rect 5122 17145 5150 19485
rect 5794 17737 5822 18773
rect 4162 17043 4286 17071
rect 5026 17117 5150 17145
rect 5698 17709 5822 17737
rect 3970 16331 3998 16923
rect 4162 16331 4190 17043
rect 3298 16229 3422 16257
rect 3682 16303 3998 16331
rect 4066 16303 4190 16331
rect 3298 15193 3326 16229
rect 3490 12973 3518 15665
rect 3682 15637 3710 16303
rect 4066 15785 4094 16303
rect 4930 15665 4958 16997
rect 5026 16969 5054 17117
rect 5698 16923 5726 17709
rect 5986 17191 6014 19069
rect 6178 18477 6206 19439
rect 7810 19041 7838 19661
rect 7426 18523 7454 18921
rect 6178 18449 6302 18477
rect 6274 17589 6302 18449
rect 6178 17561 6302 17589
rect 6178 17413 6206 17561
rect 6850 16969 6878 17741
rect 7618 17737 7646 18995
rect 7522 17709 7646 17737
rect 7522 17219 7550 17709
rect 7522 17191 7646 17219
rect 5698 16895 5822 16923
rect 5794 16775 5822 16895
rect 5794 16747 5918 16775
rect 5794 16525 5822 16747
rect 7618 16525 7646 17191
rect 7810 16493 7838 18921
rect 6082 15761 6110 16331
rect 6850 15813 6878 16331
rect 6754 15785 6878 15813
rect 3586 15517 3614 15591
rect 4258 15221 4286 15665
rect 4930 15637 5150 15665
rect 4258 15193 4574 15221
rect 3682 14994 3710 15073
rect 3682 14175 3710 14259
rect 3586 13662 3614 13741
rect 3586 12899 3614 12983
rect 3202 12307 3518 12335
rect 3010 12159 3134 12187
rect 2818 12085 2942 12113
rect 2242 11937 2366 11965
rect 2050 11641 2174 11669
rect 2050 11003 2078 11641
rect 1954 10975 2078 11003
rect 1954 10411 1982 10975
rect 2146 10457 2174 10929
rect 1954 10383 2078 10411
rect 1954 9643 1982 10115
rect 1282 9495 1406 9523
rect 1378 9005 1406 9495
rect 1282 8977 1406 9005
rect 1090 8903 1214 8931
rect 322 8533 446 8561
rect 34 8117 62 8191
rect 0 8089 97 8117
rect 226 7673 254 8265
rect 418 7673 446 8533
rect 802 8533 926 8561
rect 802 8089 830 8533
rect 0 7645 254 7673
rect 322 7645 446 7673
rect 0 7127 97 7155
rect 34 6933 62 7127
rect 34 6905 158 6933
rect 226 6785 254 7451
rect 322 6979 350 7645
rect 994 7155 1022 8783
rect 898 7127 1022 7155
rect 34 6757 254 6785
rect 34 6711 62 6757
rect 0 6683 97 6711
rect 34 6267 62 6517
rect 0 6239 97 6267
rect 34 5749 62 6193
rect 322 5749 350 6341
rect 898 6193 926 7127
rect 898 6165 1022 6193
rect 0 5721 97 5749
rect 322 5721 542 5749
rect 130 5527 158 5675
rect 34 5305 62 5527
rect 130 5499 206 5527
rect 0 5277 97 5305
rect 34 4787 62 4861
rect 0 4759 97 4787
rect 0 4315 97 4343
rect 178 4269 206 5499
rect 514 4861 542 5721
rect 322 4833 542 4861
rect 322 4491 350 4833
rect 994 4537 1022 6165
rect 1186 5869 1214 8903
rect 1282 8829 1310 8977
rect 1378 8117 1406 8265
rect 1378 8089 1502 8117
rect 1474 6933 1502 8089
rect 1762 7201 1790 8413
rect 1378 6905 1502 6933
rect 1378 6535 1406 6905
rect 1570 6415 1598 6785
rect 1474 6387 1598 6415
rect 1474 5823 1502 6387
rect 1474 5795 1598 5823
rect 1570 5647 1598 5795
rect 322 4463 542 4491
rect 130 4241 206 4269
rect 130 3899 158 4241
rect 130 3871 206 3899
rect 0 3797 97 3825
rect 0 3353 97 3381
rect 178 3307 206 3871
rect 514 3529 542 4463
rect 130 3279 206 3307
rect 322 3501 542 3529
rect 130 2937 158 3279
rect 322 3159 350 3501
rect 322 3131 446 3159
rect 130 2909 206 2937
rect 0 2835 97 2863
rect 34 2419 62 2493
rect 0 2391 97 2419
rect 34 1901 62 2197
rect 178 1975 206 2909
rect 418 2641 446 3131
rect 322 2613 446 2641
rect 322 2465 350 2613
rect 130 1947 206 1975
rect 0 1873 97 1901
rect 130 1827 158 1947
rect 34 1799 158 1827
rect 34 1457 62 1799
rect 0 1429 97 1457
rect 898 1309 926 4343
rect 1282 2983 1310 3603
rect 994 2391 1022 2789
rect 1090 1651 1118 2123
rect 34 1281 926 1309
rect 34 939 62 1281
rect 0 911 97 939
rect 34 495 62 865
rect 0 467 97 495
rect 130 421 158 1013
rect 1762 837 1790 7007
rect 2050 6313 2078 8561
rect 2338 8265 2366 11937
rect 2914 11641 2942 12085
rect 3106 11595 3134 12159
rect 3010 11567 3134 11595
rect 3010 10855 3038 11567
rect 3298 10975 3326 12187
rect 3490 11003 3518 12307
rect 4066 11743 4094 14555
rect 4546 14305 4574 15193
rect 4930 12381 4958 14333
rect 5122 13667 5150 14999
rect 5986 14379 6014 15665
rect 6754 15637 6782 15785
rect 7042 15637 7070 16331
rect 8098 15761 8126 20646
rect 8290 17811 8318 18403
rect 8290 17783 8414 17811
rect 8386 17293 8414 17783
rect 8290 17265 8414 17293
rect 8290 17103 8318 17265
rect 8290 16525 8318 16997
rect 8866 16303 8894 16997
rect 8578 15785 8606 16183
rect 6274 14259 6302 14999
rect 8098 14994 8126 15073
rect 6178 14231 6302 14259
rect 5122 13639 5246 13667
rect 5122 12973 5150 13639
rect 5986 12529 6014 13445
rect 4546 11789 4574 12261
rect 3970 11715 4094 11743
rect 3970 11151 3998 11715
rect 4258 11225 4286 11669
rect 4738 11521 4766 11669
rect 5314 11641 5342 12409
rect 5602 11567 5630 12335
rect 6178 11789 6206 14231
rect 6658 12922 6686 13001
rect 6850 11817 6878 14333
rect 7138 13639 7166 14333
rect 8098 14231 8126 14325
rect 8098 13662 8126 13741
rect 8098 12899 8126 12983
rect 8290 12973 8318 15665
rect 8962 12973 8990 15665
rect 9250 13149 9278 18329
rect 9634 16969 9662 20401
rect 12130 20373 12158 20646
rect 13378 19855 13406 20646
rect 10306 17071 10334 18773
rect 10210 17043 10334 17071
rect 10210 16035 10238 17043
rect 11362 16997 11390 18773
rect 11650 17191 11678 18847
rect 10498 16109 10526 16997
rect 11362 16969 11582 16997
rect 11362 16525 11390 16969
rect 13090 16525 13118 18773
rect 13282 18033 13310 19143
rect 13474 18995 13502 19661
rect 13474 18967 13598 18995
rect 13570 18329 13598 18967
rect 13474 18301 13598 18329
rect 13474 18153 13502 18301
rect 13282 18005 13406 18033
rect 13378 16479 13406 18005
rect 15106 17589 15134 20646
rect 17506 19855 17534 20646
rect 16834 19217 16862 19587
rect 16642 19189 16862 19217
rect 16066 18181 16094 18351
rect 15970 18153 16094 18181
rect 15490 17663 15518 18107
rect 15490 17635 15614 17663
rect 15106 17561 15326 17589
rect 10498 16081 10910 16109
rect 10210 16007 10334 16035
rect 9634 13519 9662 15221
rect 10306 15193 10334 16007
rect 10882 15785 10910 16081
rect 10306 14305 10334 15073
rect 10498 13639 10526 14333
rect 10978 14111 11006 14259
rect 10882 14083 11006 14111
rect 9154 13121 9278 13149
rect 9538 13491 9662 13519
rect 10882 13519 10910 14083
rect 11170 13593 11198 15789
rect 11650 15637 11678 16479
rect 13282 16451 13406 16479
rect 11842 14231 11870 15665
rect 12226 14971 12254 16331
rect 13282 15739 13310 16451
rect 13186 15711 13310 15739
rect 13186 15221 13214 15711
rect 13186 15193 13310 15221
rect 13090 14971 13118 15057
rect 11170 13565 11294 13593
rect 10882 13491 11006 13519
rect 9154 13001 9182 13121
rect 9058 12973 9182 13001
rect 9058 12927 9086 12973
rect 8962 12899 9086 12927
rect 6754 11789 6878 11817
rect 4738 11493 4862 11521
rect 4258 11197 4478 11225
rect 3970 11123 4094 11151
rect 3490 10975 3710 11003
rect 2962 10827 3038 10855
rect 2818 10263 2846 10411
rect 2962 10337 2990 10827
rect 3106 10383 3134 10781
rect 2962 10309 3038 10337
rect 2722 10235 2846 10263
rect 2722 9523 2750 10235
rect 2722 9495 2942 9523
rect 2914 9227 2942 9495
rect 2818 9199 2942 9227
rect 2818 8533 2846 9199
rect 2242 8237 2366 8265
rect 2242 7719 2270 8117
rect 1858 2539 1886 2937
rect 1858 1873 1886 2345
rect 1954 1651 1982 2789
rect 2050 2539 2078 3751
rect 1858 1207 1886 1605
rect 2146 1207 2174 2271
rect 2338 1059 2366 1457
rect 34 393 158 421
rect 34 51 62 393
rect 994 319 1022 791
rect 2626 393 2654 1013
rect 2914 393 2942 2123
rect 1762 267 1790 347
rect 3010 319 3038 10309
rect 3298 9791 3326 10855
rect 3490 9717 3518 10929
rect 3682 10855 3710 10975
rect 3682 10827 3806 10855
rect 3298 7155 3326 9523
rect 3490 8385 3518 9597
rect 3778 9375 3806 10827
rect 3682 9347 3806 9375
rect 3682 9199 3710 9347
rect 4066 9079 4094 11123
rect 4450 10337 4478 11197
rect 4834 10975 4862 11493
rect 6082 10975 6110 11669
rect 6370 10975 6398 11669
rect 6754 11077 6782 11789
rect 7042 11197 7070 12335
rect 6754 11049 6878 11077
rect 4354 10309 4478 10337
rect 5218 9643 5246 10337
rect 3970 9051 4094 9079
rect 3490 7303 3518 8191
rect 3490 7275 3614 7303
rect 3298 7127 3518 7155
rect 3490 5721 3518 7127
rect 3586 6979 3614 7275
rect 3970 6119 3998 9051
rect 5986 9005 6014 10909
rect 6850 10881 6878 11049
rect 7042 10383 7070 11003
rect 6466 9643 6494 10337
rect 4258 6165 4286 9005
rect 5410 8977 6014 9005
rect 3970 6091 4094 6119
rect 4066 4389 4094 6091
rect 5410 4833 5438 8977
rect 5986 5499 6014 8339
rect 6466 8117 6494 9079
rect 6274 8089 6494 8117
rect 6274 7645 6302 8089
rect 7618 6489 7646 9597
rect 7906 6979 7934 9523
rect 8098 9417 8126 9671
rect 8290 8385 8318 11669
rect 8962 11641 8990 12899
rect 9538 11595 9566 13491
rect 9826 11641 9854 13445
rect 8866 11003 8894 11595
rect 9538 11567 9662 11595
rect 8866 10975 9182 11003
rect 8866 10309 8894 10975
rect 9058 9417 9086 9671
rect 8098 7587 8126 7673
rect 9154 6979 9182 7599
rect 3106 393 3134 2419
rect 3202 393 3230 1457
rect 3874 1207 3902 1605
rect 3394 541 3422 939
rect 3778 319 3806 939
rect 9634 569 9662 11567
rect 10978 10235 11006 13491
rect 11266 10411 11294 13565
rect 11746 11641 11774 13715
rect 12130 12307 12158 13667
rect 12322 10975 12350 11743
rect 13282 11669 13310 15193
rect 13474 14999 13502 15665
rect 13666 15637 13694 16331
rect 13474 14971 13694 14999
rect 13666 12973 13694 14971
rect 13858 14333 13886 17441
rect 14338 15665 14366 17441
rect 15010 17367 15038 17497
rect 15010 17339 15134 17367
rect 15106 17145 15134 17339
rect 15010 17117 15134 17145
rect 15010 16183 15038 17117
rect 15298 16183 15326 17561
rect 15586 17145 15614 17635
rect 15490 17117 15614 17145
rect 15970 17145 15998 18153
rect 15970 17117 16094 17145
rect 15010 16155 15134 16183
rect 15298 16155 15422 16183
rect 14242 15637 14366 15665
rect 14242 14999 14270 15637
rect 14242 14971 14366 14999
rect 14530 14971 14558 15665
rect 15106 15073 15134 16155
rect 15394 16035 15422 16155
rect 15298 16007 15422 16035
rect 15298 15883 15326 16007
rect 15106 15045 15230 15073
rect 13858 14305 13982 14333
rect 13954 13667 13982 14305
rect 13858 13639 13982 13667
rect 13282 11641 13406 11669
rect 13090 10855 13118 11595
rect 11170 10383 11294 10411
rect 12994 10827 13118 10855
rect 11170 10041 11198 10383
rect 10978 10013 11198 10041
rect 10306 8977 10334 9745
rect 9634 541 9758 569
rect 5890 319 6110 347
rect 0 23 97 51
rect 5890 0 5918 319
rect 10978 0 11006 10013
rect 11362 9643 11390 10263
rect 11650 9643 11678 10337
rect 12994 9717 13022 10827
rect 13378 10781 13406 11641
rect 13858 11077 13886 13639
rect 14146 11123 14174 12261
rect 14338 11817 14366 14971
rect 14914 14555 14942 14999
rect 14626 14527 14942 14555
rect 14626 13519 14654 14527
rect 15202 14481 15230 15045
rect 15106 14453 15230 14481
rect 14626 13491 14942 13519
rect 14914 13223 14942 13491
rect 14626 13195 14942 13223
rect 14626 12335 14654 13195
rect 15106 12409 15134 14453
rect 15106 12381 15230 12409
rect 14626 12307 14942 12335
rect 14338 11789 14462 11817
rect 14434 11077 14462 11789
rect 14914 11641 14942 12307
rect 15202 11595 15230 12381
rect 13282 10753 13406 10781
rect 13762 11049 13886 11077
rect 14338 11049 14462 11077
rect 15106 11567 15230 11595
rect 11746 0 11774 4269
rect 12610 0 12638 569
rect 13282 62 13310 10753
rect 13762 10263 13790 11049
rect 14050 10309 14078 11003
rect 13762 10235 13886 10263
rect 13858 1651 13886 10235
rect 13954 1207 13982 1679
rect 14242 1059 14270 1457
rect 13378 541 13406 1013
rect 13474 62 13502 97
rect 13282 34 13502 62
rect 13474 0 13502 34
rect 14242 0 14270 199
rect 14338 171 14366 11049
rect 15106 0 15134 11567
rect 15490 2243 15518 17117
rect 15778 7571 15806 16997
rect 16066 5083 16094 17117
rect 16258 16525 16286 18847
rect 16642 18153 16670 19189
rect 17794 18893 17918 18921
rect 16450 17117 16478 17811
rect 17218 17145 17246 18107
rect 17602 17857 17630 18181
rect 17218 17117 17342 17145
rect 17026 16377 17054 17071
rect 17314 16331 17342 17117
rect 17794 17071 17822 18893
rect 19330 18477 19358 20646
rect 19618 18893 19646 20253
rect 21730 19855 21758 20646
rect 20290 19217 20318 19661
rect 20290 19189 20510 19217
rect 20098 18995 20126 19143
rect 20002 18967 20126 18995
rect 20482 18995 20510 19189
rect 20482 18967 20606 18995
rect 19330 18449 19646 18477
rect 18850 17145 18878 17515
rect 18754 17117 18878 17145
rect 17794 17043 17918 17071
rect 17794 16525 17822 17043
rect 17218 16303 17342 16331
rect 15970 5055 16094 5083
rect 15298 319 15326 791
rect 15970 0 15998 5055
rect 16066 1207 16094 1679
rect 16258 1059 16286 1531
rect 16834 569 16862 15221
rect 17218 9865 17246 16303
rect 18754 16183 18782 17117
rect 17794 15489 17822 16109
rect 18082 15637 18110 16183
rect 18754 16155 18878 16183
rect 17986 13195 18014 15591
rect 18274 10855 18302 15665
rect 18658 14971 18686 15517
rect 18850 14481 18878 16155
rect 19042 15073 19070 18107
rect 18658 14453 18878 14481
rect 18994 15045 19070 15073
rect 19330 15073 19358 18107
rect 19618 16701 19646 18449
rect 20002 17811 20030 18967
rect 20290 17885 20318 18921
rect 20578 18329 20606 18967
rect 21826 18523 21854 18921
rect 22018 18847 22046 18921
rect 21922 18819 22046 18847
rect 20482 18301 20606 18329
rect 20482 18153 20510 18301
rect 20866 17885 20894 18181
rect 20290 17857 20414 17885
rect 20002 17783 20126 17811
rect 19906 17413 19934 17497
rect 19522 16673 19646 16701
rect 19522 16155 19550 16673
rect 19330 15045 19454 15073
rect 18658 13519 18686 14453
rect 18994 14037 19022 15045
rect 18946 14009 19022 14037
rect 18946 13519 18974 14009
rect 19138 13593 19166 14999
rect 19042 13565 19166 13593
rect 18658 13491 18878 13519
rect 18946 13491 19022 13519
rect 18850 13149 18878 13491
rect 18754 13121 18878 13149
rect 18754 12187 18782 13121
rect 18994 12927 19022 13491
rect 19138 12973 19166 13565
rect 19426 12927 19454 15045
rect 18994 12899 19070 12927
rect 18754 12159 18878 12187
rect 18850 11817 18878 12159
rect 18178 10827 18302 10855
rect 18754 11789 18878 11817
rect 18754 10855 18782 11789
rect 18754 10827 18878 10855
rect 16930 1873 16958 2345
rect 17410 1651 17438 2123
rect 16930 1059 16958 1457
rect 16738 541 16862 569
rect 16738 0 16766 541
rect 17602 0 17630 7599
rect 17890 125 17918 10263
rect 18178 3233 18206 10827
rect 18850 10485 18878 10827
rect 18754 10457 18878 10485
rect 18754 9523 18782 10457
rect 18754 9495 18878 9523
rect 18850 9153 18878 9495
rect 18754 9125 18878 9153
rect 18754 8191 18782 9125
rect 18754 8163 18878 8191
rect 18850 7821 18878 8163
rect 18754 7793 18878 7821
rect 18754 6859 18782 7793
rect 18754 6831 18878 6859
rect 18850 6489 18878 6831
rect 18754 6461 18878 6489
rect 18754 5527 18782 6461
rect 18754 5499 18878 5527
rect 18850 5157 18878 5499
rect 18754 5129 18878 5157
rect 18754 4195 18782 5129
rect 18754 4167 18878 4195
rect 18850 3825 18878 4167
rect 18082 3205 18206 3233
rect 18754 3797 18878 3825
rect 18082 2493 18110 3205
rect 18754 2863 18782 3797
rect 18754 2835 18878 2863
rect 18850 2493 18878 2835
rect 18082 2465 18206 2493
rect 18178 1531 18206 2465
rect 18754 2465 18878 2493
rect 18082 1503 18206 1531
rect 18082 1235 18110 1503
rect 18082 1207 18206 1235
rect 18274 1207 18302 1679
rect 18754 1531 18782 2465
rect 18754 1503 18878 1531
rect 17890 97 18110 125
rect 18082 0 18110 97
rect 18178 0 18206 1207
rect 18850 1161 18878 1503
rect 18754 1133 18878 1161
rect 18754 421 18782 1133
rect 19042 467 19070 12899
rect 19330 12899 19454 12927
rect 18754 393 18878 421
rect 18850 245 18878 393
rect 18466 0 18494 199
rect 19330 0 19358 12899
rect 19906 10041 19934 16923
rect 20098 16627 20126 17783
rect 20386 16775 20414 17857
rect 20578 17857 20894 17885
rect 20578 17191 20606 17857
rect 21730 17293 21758 17441
rect 21634 17265 21758 17293
rect 20290 16747 20414 16775
rect 20098 16599 20222 16627
rect 19906 10013 20030 10041
rect 19714 1133 19742 9893
rect 20002 911 20030 10013
rect 20194 9819 20222 16599
rect 20290 16525 20318 16747
rect 20194 9791 20318 9819
rect 20290 8857 20318 9791
rect 20194 8829 20318 8857
rect 20194 8487 20222 8829
rect 20194 8459 20318 8487
rect 20290 7525 20318 8459
rect 20194 7497 20318 7525
rect 20194 7155 20222 7497
rect 20194 7127 20318 7155
rect 20290 6193 20318 7127
rect 20194 6165 20318 6193
rect 20194 5823 20222 6165
rect 20194 5795 20318 5823
rect 20290 4861 20318 5795
rect 20194 4833 20318 4861
rect 20194 4491 20222 4833
rect 20194 4463 20318 4491
rect 20290 3529 20318 4463
rect 20194 3501 20318 3529
rect 20194 3159 20222 3501
rect 20194 3131 20318 3159
rect 20290 2197 20318 3131
rect 20194 2169 20318 2197
rect 20194 1827 20222 2169
rect 20194 1799 20318 1827
rect 20290 865 20318 1799
rect 20098 837 20318 865
rect 20098 0 20126 837
rect 20962 0 20990 16775
rect 21634 13371 21662 17265
rect 21922 16525 21950 18819
rect 22306 17191 22334 17811
rect 21634 13343 21758 13371
rect 21730 13195 21758 13343
rect 21922 10235 21950 16109
rect 22114 15591 22142 16183
rect 22306 15637 22334 16331
rect 22114 15563 22238 15591
rect 22210 14994 22238 15563
rect 22306 13223 22334 14111
rect 22306 13195 22430 13223
rect 22402 13047 22430 13195
rect 22882 11715 22910 15073
rect 22978 12973 23006 15665
rect 23266 12187 23294 14925
rect 23458 13667 23486 18773
rect 24034 14971 24062 15665
rect 24130 15193 24158 16331
rect 23170 12159 23294 12187
rect 23362 13639 23486 13667
rect 23170 11863 23198 12159
rect 23266 11715 23294 12113
rect 23362 11003 23390 13639
rect 23554 12307 23582 12853
rect 23650 11049 23678 13593
rect 23362 10975 23486 11003
rect 21730 1577 21854 1605
rect 21826 0 21854 1577
rect 22306 1235 22334 2197
rect 22306 1207 22622 1235
rect 22594 0 22622 1207
rect 23458 0 23486 10975
rect 23746 10929 23774 14777
rect 24130 13713 24158 14259
rect 24322 13815 24350 17145
rect 24514 15859 24542 16331
rect 24706 14999 24734 15147
rect 24706 14971 24830 14999
rect 24802 14333 24830 14971
rect 24994 14925 25022 15591
rect 24898 14897 25022 14925
rect 24898 14527 24926 14897
rect 24802 14305 24926 14333
rect 24322 13787 24446 13815
rect 23650 10901 23774 10929
rect 23842 10235 23870 13593
rect 24034 13519 24062 13667
rect 23986 13491 24062 13519
rect 23986 12335 24014 13491
rect 24130 12381 24158 13445
rect 24226 12529 24254 13001
rect 24418 12853 24446 13787
rect 24898 13639 24926 14305
rect 25186 13297 25214 15665
rect 25474 13713 25502 14259
rect 25186 13269 25310 13297
rect 24322 12825 24446 12853
rect 23986 12307 24062 12335
rect 24034 11567 24062 12307
rect 24130 11197 24158 12261
rect 24322 0 24350 12825
rect 24994 12483 25022 13223
rect 24898 12455 25022 12483
rect 24898 11743 24926 12455
rect 25282 12409 25310 13269
rect 25186 12381 25310 12409
rect 25186 11817 25214 12381
rect 25186 11789 25310 11817
rect 25570 11789 25598 14999
rect 25666 13047 25694 14555
rect 25762 13047 25790 14111
rect 25762 12187 25790 12335
rect 25666 12159 25790 12187
rect 24898 11715 25022 11743
rect 24994 5083 25022 11715
rect 25282 5157 25310 11789
rect 25666 11669 25694 12159
rect 25858 11863 25886 13001
rect 25666 11641 25790 11669
rect 25762 10309 25790 11641
rect 25282 5129 25406 5157
rect 24994 5055 25118 5083
rect 25090 4491 25118 5055
rect 24994 4463 25118 4491
rect 24994 3529 25022 4463
rect 25378 4417 25406 5129
rect 25282 4389 25406 4417
rect 25282 3603 25310 4389
rect 25282 3575 25406 3603
rect 24994 3501 25118 3529
rect 25090 3159 25118 3501
rect 24994 3131 25118 3159
rect 24994 2197 25022 3131
rect 25378 3085 25406 3575
rect 25282 3057 25406 3085
rect 25282 2271 25310 3057
rect 25282 2243 25406 2271
rect 24994 2169 25118 2197
rect 25090 1827 25118 2169
rect 24994 1799 25118 1827
rect 24994 865 25022 1799
rect 25378 1753 25406 2243
rect 25282 1725 25406 1753
rect 24994 837 25118 865
rect 25090 0 25118 837
rect 25282 393 25310 1725
rect 25954 0 25982 18329
rect 26914 15665 26942 18551
rect 26818 15637 26942 15665
rect 26818 14851 26846 15637
rect 26818 14823 26942 14851
rect 27106 14823 27134 15591
rect 26626 13861 26654 14333
rect 26146 11641 26174 12113
rect 26146 10975 26174 11447
rect 26242 10975 26270 12927
rect 26146 10457 26174 10781
rect 26914 1235 26942 14823
rect 27010 12529 27038 14185
rect 27202 13713 27230 14777
rect 27394 14231 27422 14925
rect 27394 12455 27422 12779
rect 27682 12187 27710 16997
rect 28066 15295 28094 15443
rect 27970 15267 28094 15295
rect 27970 12335 27998 15267
rect 28258 12409 28286 17441
rect 28258 12381 28382 12409
rect 27970 12307 28094 12335
rect 27682 12159 27806 12187
rect 27490 11641 27518 12113
rect 27010 11197 27038 11595
rect 27490 10975 27518 11447
rect 27490 10309 27518 10781
rect 27778 10263 27806 12159
rect 26818 1207 26942 1235
rect 27682 10235 27806 10263
rect 26818 0 26846 1207
rect 27682 0 27710 10235
rect 28066 9783 28094 12307
rect 28354 11521 28382 12381
rect 28642 11715 28670 12261
rect 28258 11493 28382 11521
rect 28258 11151 28286 11493
rect 28258 11123 28382 11151
rect 28354 10189 28382 11123
rect 28834 11049 28862 12113
rect 29026 10235 29054 15665
rect 28258 10161 28382 10189
rect 28258 569 28286 10161
rect 28258 541 28478 569
rect 28450 0 28478 541
rect 29314 0 29342 18255
rect 29794 14971 29822 15443
rect 29890 14305 29918 14777
rect 29698 13639 29726 14111
rect 29794 13593 29822 13741
rect 29698 13565 29822 13593
rect 29602 12233 29630 12927
rect 29698 10975 29726 13565
rect 30178 0 30206 18773
rect 30946 0 30974 16331
rect 32866 569 32894 1087
rect 32674 541 32894 569
rect 31810 0 31838 199
rect 32674 0 32702 541
rect 33442 0 33470 18921
rect 34018 837 34334 865
rect 34306 0 34334 837
rect 35170 0 35198 17253
rect 35938 0 35966 495
<< metal3 >>
rect 18 19771 5070 19831
rect 18 18795 4590 18855
rect 4146 18307 16110 18367
rect 18 17819 270 17879
rect 210 17757 270 17819
rect 5010 17819 6606 17879
rect 5010 17757 5070 17819
rect 210 17697 5070 17757
rect 6546 17757 6606 17819
rect 6546 17697 6894 17757
rect 4434 17453 15054 17513
rect 19890 17453 35214 17513
rect 35154 17209 35214 17453
rect 18 17087 8334 17147
rect 3762 16843 8334 16903
rect 18 16477 7854 16537
rect 1266 16111 11214 16171
rect 6066 15745 8142 15805
rect 11154 15745 11214 16111
rect 15282 15867 17934 15927
rect 3473 15501 3630 15561
rect 3522 15013 3726 15073
rect 7990 15013 8112 15073
rect 13074 15013 14142 15073
rect 22102 15013 22224 15073
rect 498 14281 1710 14341
rect 7990 14281 8112 14341
rect 978 13731 1038 14281
rect 3522 14159 3726 14219
rect 17873 14159 18030 14219
rect 498 13671 1038 13731
rect 3473 13671 3630 13731
rect 7990 13671 8112 13731
rect 10482 13671 11790 13731
rect 22194 13061 22446 13121
rect 3473 12939 3630 12999
rect 5970 12939 6702 12999
rect 7990 12939 8112 12999
rect 12114 12817 14142 12877
rect 18 12329 1902 12389
rect 1510 11597 1662 11657
rect 1170 11109 6126 11169
rect 5970 10865 6894 10925
rect 14034 10865 17934 10925
rect 978 10255 1230 10315
rect 978 10193 1038 10255
rect 18 10133 1038 10193
rect 978 10071 1038 10133
rect 978 10011 1230 10071
rect 1170 9827 1230 10011
rect 1170 9767 28110 9827
rect 7990 9401 9102 9461
rect 7990 7571 8112 7631
rect 18 6473 7662 6533
rect 1602 251 1806 311
<< metal4 >>
rect 1602 251 1662 11657
rect 3452 6660 3652 15984
rect 7964 6660 8164 15984
rect 14012 6660 14212 15984
rect 17852 6660 18052 15984
rect 22076 6660 22276 15984
<< metal5 >>
rect 400 0 800 20646
rect 2400 0 2800 20646
rect 4400 0 4800 20646
rect 6400 0 6800 20646
rect 8400 0 8800 20646
rect 10400 0 10800 20646
rect 12400 0 12800 20646
rect 14400 0 14800 20646
rect 16400 0 16800 20646
rect 18400 0 18800 20646
rect 20400 0 20800 20646
rect 22400 0 22800 20646
rect 24400 0 24800 20646
rect 26400 0 26800 20646
rect 28400 0 28800 20646
rect 30400 0 30800 20646
rect 32400 0 32800 20646
rect 34400 0 34800 20646
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_258
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_517
timestamp 1626908933
transform 1 0 288 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_256
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_624
timestamp 1626908933
transform 1 0 384 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_441
timestamp 1626908933
transform 1 0 576 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1071
timestamp 1626908933
transform 1 0 576 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_4
timestamp 1626908933
transform 1 0 672 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_44
timestamp 1626908933
transform 1 0 672 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_41
timestamp 1626908933
transform 1 0 1440 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_1
timestamp 1626908933
transform 1 0 1440 0 1 0
box -38 -49 806 715
use M3M4_PR  M3M4_PR_41
timestamp 1626908933
transform 1 0 1632 0 1 281
box -38 -33 38 33
use M3M4_PR  M3M4_PR_20
timestamp 1626908933
transform 1 0 1632 0 1 281
box -38 -33 38 33
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1070
timestamp 1626908933
transform 1 0 2208 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_440
timestamp 1626908933
transform 1 0 2208 0 1 0
box -38 -49 134 715
use M2M3_PR  M2M3_PR_86
timestamp 1626908933
transform 1 0 1776 0 1 281
box -33 -37 33 37
use M2M3_PR  M2M3_PR_27
timestamp 1626908933
transform 1 0 1776 0 1 281
box -33 -37 33 37
use osc_core_VIA10  osc_core_VIA10_27
timestamp 1626908933
transform 1 0 2600 0 1 23
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_13
timestamp 1626908933
transform 1 0 2600 0 1 23
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_27
timestamp 1626908933
transform 1 0 2600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_13
timestamp 1626908933
transform 1 0 2600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_35
timestamp 1626908933
transform 1 0 2600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_17
timestamp 1626908933
transform 1 0 2600 0 1 16
box -200 -33 200 33
use osc_core_VIA4  osc_core_VIA4_287
timestamp 1626908933
transform 1 0 2600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_575
timestamp 1626908933
transform 1 0 2600 0 1 93
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_516
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_257
timestamp 1626908933
transform 1 0 2496 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_625
timestamp 1626908933
transform 1 0 2304 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_257
timestamp 1626908933
transform 1 0 2304 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_14
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_5
timestamp 1626908933
transform 1 0 2592 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_15
timestamp 1626908933
transform 1 0 2976 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_6
timestamp 1626908933
transform 1 0 2976 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__buf_4  sky130_fd_sc_hs__buf_4_0
timestamp 1626908933
transform 1 0 3360 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__buf_4  sky130_fd_sc_hs__buf_4_1
timestamp 1626908933
transform 1 0 3360 0 1 0
box -38 -49 710 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1114
timestamp 1626908933
transform 1 0 4032 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_544
timestamp 1626908933
transform 1 0 4032 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_515
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_256
timestamp 1626908933
transform 1 0 4992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1072
timestamp 1626908933
transform 1 0 4896 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1060
timestamp 1626908933
transform 1 0 4800 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_442
timestamp 1626908933
transform 1 0 4896 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_430
timestamp 1626908933
transform 1 0 4800 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1100
timestamp 1626908933
transform 1 0 5280 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_530
timestamp 1626908933
transform 1 0 5280 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_621
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_253
timestamp 1626908933
transform 1 0 5088 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_429
timestamp 1626908933
transform 1 0 6048 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1059
timestamp 1626908933
transform 1 0 6048 0 1 0
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_559
timestamp 1626908933
transform 1 0 6600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_271
timestamp 1626908933
transform 1 0 6600 0 1 93
box -200 -142 200 178
use osc_core_VIA10  osc_core_VIA10_26
timestamp 1626908933
transform 1 0 6600 0 1 23
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_12
timestamp 1626908933
transform 1 0 6600 0 1 23
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_26
timestamp 1626908933
transform 1 0 6600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_12
timestamp 1626908933
transform 1 0 6600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_34
timestamp 1626908933
transform 1 0 6600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_16
timestamp 1626908933
transform 1 0 6600 0 1 16
box -200 -33 200 33
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1058
timestamp 1626908933
transform 1 0 6528 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_428
timestamp 1626908933
transform 1 0 6528 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_516
timestamp 1626908933
transform 1 0 6624 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1086
timestamp 1626908933
transform 1 0 6624 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_505
timestamp 1626908933
transform 1 0 6144 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1074
timestamp 1626908933
transform 1 0 6144 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1057
timestamp 1626908933
transform 1 0 7776 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_427
timestamp 1626908933
transform 1 0 7776 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1073
timestamp 1626908933
transform 1 0 7392 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_443
timestamp 1626908933
transform 1 0 7392 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_514
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_255
timestamp 1626908933
transform 1 0 7488 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_620
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_252
timestamp 1626908933
transform 1 0 7584 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1070
timestamp 1626908933
transform 1 0 7872 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_500
timestamp 1626908933
transform 1 0 7872 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1049
timestamp 1626908933
transform 1 0 8736 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_480
timestamp 1626908933
transform 1 0 8736 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1056
timestamp 1626908933
transform 1 0 9120 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_486
timestamp 1626908933
transform 1 0 9120 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1056
timestamp 1626908933
transform 1 0 8640 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_426
timestamp 1626908933
transform 1 0 8640 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_254
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_513
timestamp 1626908933
transform 1 0 9984 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_444
timestamp 1626908933
transform 1 0 9888 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1074
timestamp 1626908933
transform 1 0 9888 0 1 0
box -38 -49 134 715
use osc_core_VIA8  osc_core_VIA8_15
timestamp 1626908933
transform 1 0 10600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_33
timestamp 1626908933
transform 1 0 10600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_11
timestamp 1626908933
transform 1 0 10600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_25
timestamp 1626908933
transform 1 0 10600 0 1 16
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_11
timestamp 1626908933
transform 1 0 10600 0 1 23
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_25
timestamp 1626908933
transform 1 0 10600 0 1 23
box -200 -26 200 26
use osc_core_VIA4  osc_core_VIA4_255
timestamp 1626908933
transform 1 0 10600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_543
timestamp 1626908933
transform 1 0 10600 0 1 93
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_473
timestamp 1626908933
transform 1 0 10464 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1043
timestamp 1626908933
transform 1 0 10464 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_453
timestamp 1626908933
transform 1 0 10080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1022
timestamp 1626908933
transform 1 0 10080 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1004
timestamp 1626908933
transform 1 0 11328 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_435
timestamp 1626908933
transform 1 0 11328 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1055
timestamp 1626908933
transform 1 0 11232 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_425
timestamp 1626908933
transform 1 0 11232 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1022
timestamp 1626908933
transform 1 0 11712 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_452
timestamp 1626908933
transform 1 0 11712 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_58
timestamp 1626908933
transform 1 0 12672 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_18
timestamp 1626908933
transform 1 0 12672 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1069
timestamp 1626908933
transform 1 0 12576 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_439
timestamp 1626908933
transform 1 0 12576 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_512
timestamp 1626908933
transform 1 0 12480 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_253
timestamp 1626908933
transform 1 0 12480 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_55
timestamp 1626908933
transform 1 0 13440 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_15
timestamp 1626908933
transform 1 0 13440 0 1 0
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_239
timestamp 1626908933
transform 1 0 14600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_527
timestamp 1626908933
transform 1 0 14600 0 1 93
box -200 -142 200 178
use osc_core_VIA10  osc_core_VIA10_24
timestamp 1626908933
transform 1 0 14600 0 1 23
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_10
timestamp 1626908933
transform 1 0 14600 0 1 23
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_24
timestamp 1626908933
transform 1 0 14600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_10
timestamp 1626908933
transform 1 0 14600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_32
timestamp 1626908933
transform 1 0 14600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_14
timestamp 1626908933
transform 1 0 14600 0 1 16
box -200 -33 200 33
use M1M2_PR  M1M2_PR_1338
timestamp 1626908933
transform 1 0 14256 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_570
timestamp 1626908933
transform 1 0 14256 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1351
timestamp 1626908933
transform 1 0 14352 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_583
timestamp 1626908933
transform 1 0 14352 0 1 185
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_252
timestamp 1626908933
transform 1 0 14976 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_511
timestamp 1626908933
transform 1 0 14976 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_12
timestamp 1626908933
transform 1 0 14208 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_52
timestamp 1626908933
transform 1 0 14208 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_974
timestamp 1626908933
transform 1 0 15072 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_404
timestamp 1626908933
transform 1 0 15072 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_49
timestamp 1626908933
transform 1 0 15840 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_9
timestamp 1626908933
transform 1 0 15840 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_946
timestamp 1626908933
transform 1 0 16704 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_376
timestamp 1626908933
transform 1 0 16704 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1054
timestamp 1626908933
transform 1 0 16608 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_424
timestamp 1626908933
transform 1 0 16608 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_510
timestamp 1626908933
transform 1 0 17472 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_251
timestamp 1626908933
transform 1 0 17472 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_885
timestamp 1626908933
transform 1 0 17760 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_316
timestamp 1626908933
transform 1 0 17760 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_619
timestamp 1626908933
transform 1 0 17568 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_251
timestamp 1626908933
transform 1 0 17568 0 1 0
box -38 -49 230 715
use osc_core_VIA8  osc_core_VIA8_13
timestamp 1626908933
transform 1 0 18600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_31
timestamp 1626908933
transform 1 0 18600 0 1 16
box -200 -33 200 33
use osc_core_VIA11  osc_core_VIA11_0
timestamp 1626908933
transform 1 0 18661 0 1 16
box -139 -33 139 33
use osc_core_VIA11  osc_core_VIA11_1
timestamp 1626908933
transform 1 0 18661 0 1 16
box -139 -33 139 33
use osc_core_VIA12  osc_core_VIA12_0
timestamp 1626908933
transform 1 0 18661 0 1 23
box -139 -26 139 26
use osc_core_VIA12  osc_core_VIA12_1
timestamp 1626908933
transform 1 0 18661 0 1 23
box -139 -26 139 26
use M1M2_PR  M1M2_PR_581
timestamp 1626908933
transform 1 0 18480 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1349
timestamp 1626908933
transform 1 0 18480 0 1 185
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_223
timestamp 1626908933
transform 1 0 18600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_511
timestamp 1626908933
transform 1 0 18600 0 1 93
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_354
timestamp 1626908933
transform 1 0 18144 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_924
timestamp 1626908933
transform 1 0 18144 0 1 0
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1379
timestamp 1626908933
transform 1 0 18864 0 1 259
box -32 -32 32 32
use M1M2_PR  M1M2_PR_611
timestamp 1626908933
transform 1 0 18864 0 1 259
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1068
timestamp 1626908933
transform 1 0 19104 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_438
timestamp 1626908933
transform 1 0 19104 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_618
timestamp 1626908933
transform 1 0 18912 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_250
timestamp 1626908933
transform 1 0 18912 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_46
timestamp 1626908933
transform 1 0 19200 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_6
timestamp 1626908933
transform 1 0 19200 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_623
timestamp 1626908933
transform 1 0 20064 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_255
timestamp 1626908933
transform 1 0 20064 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_509
timestamp 1626908933
transform 1 0 19968 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_250
timestamp 1626908933
transform 1 0 19968 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_43
timestamp 1626908933
transform 1 0 20256 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_3
timestamp 1626908933
transform 1 0 20256 0 1 0
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1309
timestamp 1626908933
transform 1 0 20304 0 1 259
box -29 -23 29 23
use L1M1_PR  L1M1_PR_521
timestamp 1626908933
transform 1 0 20304 0 1 259
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1053
timestamp 1626908933
transform 1 0 21024 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_423
timestamp 1626908933
transform 1 0 21024 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_831
timestamp 1626908933
transform 1 0 21120 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_262
timestamp 1626908933
transform 1 0 21120 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1067
timestamp 1626908933
transform 1 0 21600 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_437
timestamp 1626908933
transform 1 0 21600 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1052
timestamp 1626908933
transform 1 0 21504 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_422
timestamp 1626908933
transform 1 0 21504 0 1 0
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1305
timestamp 1626908933
transform 1 0 21744 0 1 259
box -29 -23 29 23
use L1M1_PR  L1M1_PR_517
timestamp 1626908933
transform 1 0 21744 0 1 259
box -29 -23 29 23
use osc_core_VIA14  osc_core_VIA14_1
timestamp 1626908933
transform 1 0 22483 0 1 23
box -83 -26 83 26
use osc_core_VIA14  osc_core_VIA14_0
timestamp 1626908933
transform 1 0 22483 0 1 23
box -83 -26 83 26
use osc_core_VIA13  osc_core_VIA13_1
timestamp 1626908933
transform 1 0 22483 0 1 16
box -83 -33 83 33
use osc_core_VIA13  osc_core_VIA13_0
timestamp 1626908933
transform 1 0 22483 0 1 16
box -83 -33 83 33
use osc_core_VIA4  osc_core_VIA4_495
timestamp 1626908933
transform 1 0 22600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_207
timestamp 1626908933
transform 1 0 22600 0 1 93
box -200 -142 200 178
use osc_core_VIA8  osc_core_VIA8_30
timestamp 1626908933
transform 1 0 22600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_12
timestamp 1626908933
transform 1 0 22600 0 1 16
box -200 -33 200 33
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_0
timestamp 1626908933
transform 1 0 21696 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_40
timestamp 1626908933
transform 1 0 21696 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_834
timestamp 1626908933
transform 1 0 22656 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_264
timestamp 1626908933
transform 1 0 22656 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1051
timestamp 1626908933
transform 1 0 22560 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_421
timestamp 1626908933
transform 1 0 22560 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_508
timestamp 1626908933
transform 1 0 22464 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_249
timestamp 1626908933
transform 1 0 22464 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_799
timestamp 1626908933
transform 1 0 23424 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_230
timestamp 1626908933
transform 1 0 23424 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1050
timestamp 1626908933
transform 1 0 23808 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_420
timestamp 1626908933
transform 1 0 23808 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_811
timestamp 1626908933
transform 1 0 23904 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_241
timestamp 1626908933
transform 1 0 23904 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_616
timestamp 1626908933
transform 1 0 25056 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_248
timestamp 1626908933
transform 1 0 25056 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_507
timestamp 1626908933
transform 1 0 24960 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_248
timestamp 1626908933
transform 1 0 24960 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_617
timestamp 1626908933
transform 1 0 24672 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_249
timestamp 1626908933
transform 1 0 24672 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1075
timestamp 1626908933
transform 1 0 24864 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_445
timestamp 1626908933
transform 1 0 24864 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_790
timestamp 1626908933
transform 1 0 25248 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_220
timestamp 1626908933
transform 1 0 25248 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_762
timestamp 1626908933
transform 1 0 26016 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_193
timestamp 1626908933
transform 1 0 26016 0 1 0
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_479
timestamp 1626908933
transform 1 0 26600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_191
timestamp 1626908933
transform 1 0 26600 0 1 93
box -200 -142 200 178
use osc_core_VIA16  osc_core_VIA16_1
timestamp 1626908933
transform 1 0 26595 0 1 23
box -195 -26 195 26
use osc_core_VIA16  osc_core_VIA16_0
timestamp 1626908933
transform 1 0 26595 0 1 23
box -195 -26 195 26
use osc_core_VIA15  osc_core_VIA15_1
timestamp 1626908933
transform 1 0 26595 0 1 16
box -195 -33 195 33
use osc_core_VIA15  osc_core_VIA15_0
timestamp 1626908933
transform 1 0 26595 0 1 16
box -195 -33 195 33
use osc_core_VIA8  osc_core_VIA8_29
timestamp 1626908933
transform 1 0 26600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_11
timestamp 1626908933
transform 1 0 26600 0 1 16
box -200 -33 200 33
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1049
timestamp 1626908933
transform 1 0 26400 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_419
timestamp 1626908933
transform 1 0 26400 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_198
timestamp 1626908933
transform 1 0 26496 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_768
timestamp 1626908933
transform 1 0 26496 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_247
timestamp 1626908933
transform 1 0 27552 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_615
timestamp 1626908933
transform 1 0 27552 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_418
timestamp 1626908933
transform 1 0 27264 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1048
timestamp 1626908933
transform 1 0 27264 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_247
timestamp 1626908933
transform 1 0 27456 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_506
timestamp 1626908933
transform 1 0 27456 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_446
timestamp 1626908933
transform 1 0 27360 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1076
timestamp 1626908933
transform 1 0 27360 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_417
timestamp 1626908933
transform 1 0 27744 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1047
timestamp 1626908933
transform 1 0 27744 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_176
timestamp 1626908933
transform 1 0 27840 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_746
timestamp 1626908933
transform 1 0 27840 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_725
timestamp 1626908933
transform 1 0 28608 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_156
timestamp 1626908933
transform 1 0 28608 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1046
timestamp 1626908933
transform 1 0 28992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_416
timestamp 1626908933
transform 1 0 28992 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_722
timestamp 1626908933
transform 1 0 29088 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_152
timestamp 1626908933
transform 1 0 29088 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1077
timestamp 1626908933
transform 1 0 29856 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_447
timestamp 1626908933
transform 1 0 29856 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_415
timestamp 1626908933
transform 1 0 30240 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1045
timestamp 1626908933
transform 1 0 30240 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_246
timestamp 1626908933
transform 1 0 29952 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_505
timestamp 1626908933
transform 1 0 29952 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_246
timestamp 1626908933
transform 1 0 30048 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_614
timestamp 1626908933
transform 1 0 30048 0 1 0
box -38 -49 230 715
use osc_core_VIA8  osc_core_VIA8_10
timestamp 1626908933
transform 1 0 30600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_28
timestamp 1626908933
transform 1 0 30600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_9
timestamp 1626908933
transform 1 0 30600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_23
timestamp 1626908933
transform 1 0 30600 0 1 16
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_9
timestamp 1626908933
transform 1 0 30600 0 1 23
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_23
timestamp 1626908933
transform 1 0 30600 0 1 23
box -200 -26 200 26
use osc_core_VIA4  osc_core_VIA4_175
timestamp 1626908933
transform 1 0 30600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_463
timestamp 1626908933
transform 1 0 30600 0 1 93
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_128
timestamp 1626908933
transform 1 0 30336 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_698
timestamp 1626908933
transform 1 0 30336 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_613
timestamp 1626908933
transform 1 0 31104 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_245
timestamp 1626908933
transform 1 0 31104 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_681
timestamp 1626908933
transform 1 0 31296 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_112
timestamp 1626908933
transform 1 0 31296 0 1 0
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1377
timestamp 1626908933
transform 1 0 31824 0 1 185
box -32 -32 32 32
use M1M2_PR  M1M2_PR_609
timestamp 1626908933
transform 1 0 31824 0 1 185
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_673
timestamp 1626908933
transform 1 0 31680 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_103
timestamp 1626908933
transform 1 0 31680 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_649
timestamp 1626908933
transform 1 0 32544 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_80
timestamp 1626908933
transform 1 0 32544 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_504
timestamp 1626908933
transform 1 0 32448 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_245
timestamp 1626908933
transform 1 0 32448 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_644
timestamp 1626908933
transform 1 0 32928 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_74
timestamp 1626908933
transform 1 0 32928 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1044
timestamp 1626908933
transform 1 0 33696 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_414
timestamp 1626908933
transform 1 0 33696 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_616
timestamp 1626908933
transform 1 0 33792 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_47
timestamp 1626908933
transform 1 0 33792 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_614
timestamp 1626908933
transform 1 0 34176 0 1 0
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_44
timestamp 1626908933
transform 1 0 34176 0 1 0
box -38 -49 806 715
use osc_core_VIA10  osc_core_VIA10_22
timestamp 1626908933
transform 1 0 34600 0 1 23
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_8
timestamp 1626908933
transform 1 0 34600 0 1 23
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_22
timestamp 1626908933
transform 1 0 34600 0 1 16
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_8
timestamp 1626908933
transform 1 0 34600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_27
timestamp 1626908933
transform 1 0 34600 0 1 16
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_9
timestamp 1626908933
transform 1 0 34600 0 1 16
box -200 -33 200 33
use osc_core_VIA4  osc_core_VIA4_159
timestamp 1626908933
transform 1 0 34600 0 1 93
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_447
timestamp 1626908933
transform 1 0 34600 0 1 93
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_244
timestamp 1626908933
transform 1 0 34944 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_503
timestamp 1626908933
transform 1 0 34944 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_258
timestamp 1626908933
transform 1 0 35424 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_626
timestamp 1626908933
transform 1 0 35424 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_448
timestamp 1626908933
transform 1 0 35616 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1078
timestamp 1626908933
transform 1 0 35616 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_15
timestamp 1626908933
transform 1 0 35040 0 1 0
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_584
timestamp 1626908933
transform 1 0 35040 0 1 0
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1535
timestamp 1626908933
transform 1 0 144 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1534
timestamp 1626908933
transform 1 0 48 0 1 851
box -32 -32 32 32
use M1M2_PR  M1M2_PR_767
timestamp 1626908933
transform 1 0 144 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_766
timestamp 1626908933
transform 1 0 48 0 1 851
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_47
timestamp 1626908933
transform 1 0 288 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_7
timestamp 1626908933
transform 1 0 288 0 -1 1332
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_134
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_404
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_134
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_404
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_134
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_404
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_143
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_431
timestamp 1626908933
transform 1 0 600 0 1 666
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1312
timestamp 1626908933
transform 1 0 816 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_524
timestamp 1626908933
transform 1 0 816 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1311
timestamp 1626908933
transform 1 0 1008 0 1 777
box -29 -23 29 23
use L1M1_PR  L1M1_PR_523
timestamp 1626908933
transform 1 0 1008 0 1 777
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1229
timestamp 1626908933
transform 1 0 1008 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_461
timestamp 1626908933
transform 1 0 1008 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1230
timestamp 1626908933
transform 1 0 1008 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_462
timestamp 1626908933
transform 1 0 1008 0 1 333
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1066
timestamp 1626908933
transform 1 0 1056 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_436
timestamp 1626908933
transform 1 0 1056 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_25
timestamp 1626908933
transform 1 0 1152 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_65
timestamp 1626908933
transform 1 0 1152 0 -1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1533
timestamp 1626908933
transform 1 0 1776 0 1 851
box -32 -32 32 32
use M1M2_PR  M1M2_PR_765
timestamp 1626908933
transform 1 0 1776 0 1 851
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1222
timestamp 1626908933
transform 1 0 1776 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_454
timestamp 1626908933
transform 1 0 1776 0 1 333
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1377
timestamp 1626908933
transform 1 0 2160 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_589
timestamp 1626908933
transform 1 0 2160 0 1 925
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_1
timestamp 1626908933
transform 1 0 1920 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_10
timestamp 1626908933
transform 1 0 1920 0 -1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1300
timestamp 1626908933
transform 1 0 2160 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_512
timestamp 1626908933
transform 1 0 2160 0 1 333
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1065
timestamp 1626908933
transform 1 0 2304 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_435
timestamp 1626908933
transform 1 0 2304 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_243
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_502
timestamp 1626908933
transform 1 0 2496 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_449
timestamp 1626908933
transform 1 0 2400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1079
timestamp 1626908933
transform 1 0 2400 0 -1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_530
timestamp 1626908933
transform 1 0 2640 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1298
timestamp 1626908933
transform 1 0 2640 0 1 407
box -32 -32 32 32
use L1M1_PR  L1M1_PR_605
timestamp 1626908933
transform 1 0 2736 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1393
timestamp 1626908933
transform 1 0 2736 0 1 407
box -29 -23 29 23
use M1M2_PR  M1M2_PR_529
timestamp 1626908933
transform 1 0 2640 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1297
timestamp 1626908933
transform 1 0 2640 0 1 999
box -32 -32 32 32
use L1M1_PR  L1M1_PR_588
timestamp 1626908933
transform 1 0 2736 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1376
timestamp 1626908933
transform 1 0 2736 0 1 925
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_11
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_2
timestamp 1626908933
transform 1 0 2592 0 -1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1300
timestamp 1626908933
transform 1 0 2928 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_532
timestamp 1626908933
transform 1 0 2928 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1302
timestamp 1626908933
transform 1 0 3120 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_534
timestamp 1626908933
transform 1 0 3120 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1340
timestamp 1626908933
transform 1 0 3024 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_572
timestamp 1626908933
transform 1 0 3024 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1304
timestamp 1626908933
transform 1 0 3216 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_536
timestamp 1626908933
transform 1 0 3216 0 1 407
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1395
timestamp 1626908933
transform 1 0 2832 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_607
timestamp 1626908933
transform 1 0 2832 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1397
timestamp 1626908933
transform 1 0 3120 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_609
timestamp 1626908933
transform 1 0 3120 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1399
timestamp 1626908933
transform 1 0 3216 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_611
timestamp 1626908933
transform 1 0 3216 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_593
timestamp 1626908933
transform 1 0 2832 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1381
timestamp 1626908933
transform 1 0 2832 0 1 925
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_535
timestamp 1626908933
transform 1 0 2976 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1104
timestamp 1626908933
transform 1 0 2976 0 -1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_520
timestamp 1626908933
transform 1 0 3408 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1288
timestamp 1626908933
transform 1 0 3408 0 1 555
box -32 -32 32 32
use L1M1_PR  L1M1_PR_592
timestamp 1626908933
transform 1 0 3504 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1380
timestamp 1626908933
transform 1 0 3504 0 1 555
box -29 -23 29 23
use M1M2_PR  M1M2_PR_519
timestamp 1626908933
transform 1 0 3408 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1287
timestamp 1626908933
transform 1 0 3408 0 1 925
box -32 -32 32 32
use L1M1_PR  L1M1_PR_601
timestamp 1626908933
transform 1 0 3504 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_604
timestamp 1626908933
transform 1 0 3600 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1389
timestamp 1626908933
transform 1 0 3504 0 1 925
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1392
timestamp 1626908933
transform 1 0 3600 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_12
timestamp 1626908933
transform 1 0 3360 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_3
timestamp 1626908933
transform 1 0 3360 0 -1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_528
timestamp 1626908933
transform 1 0 3792 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1296
timestamp 1626908933
transform 1 0 3792 0 1 333
box -32 -32 32 32
use L1M1_PR  L1M1_PR_600
timestamp 1626908933
transform 1 0 3888 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1388
timestamp 1626908933
transform 1 0 3888 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_527
timestamp 1626908933
transform 1 0 3792 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1295
timestamp 1626908933
transform 1 0 3792 0 1 925
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_413
timestamp 1626908933
transform 1 0 4128 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1043
timestamp 1626908933
transform 1 0 4128 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_17
timestamp 1626908933
transform 1 0 3744 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_8
timestamp 1626908933
transform 1 0 3744 0 -1 1332
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_119
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_389
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_119
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_389
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_119
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_389
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_127
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_415
timestamp 1626908933
transform 1 0 4600 0 1 666
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_533
timestamp 1626908933
transform 1 0 4608 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1103
timestamp 1626908933
transform 1 0 4608 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_523
timestamp 1626908933
transform 1 0 4224 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1092
timestamp 1626908933
transform 1 0 4224 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_612
timestamp 1626908933
transform 1 0 5760 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_244
timestamp 1626908933
transform 1 0 5760 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1086
timestamp 1626908933
transform 1 0 5376 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_517
timestamp 1626908933
transform 1 0 5376 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1088
timestamp 1626908933
transform 1 0 5952 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_518
timestamp 1626908933
transform 1 0 5952 0 -1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1325
timestamp 1626908933
transform 1 0 6096 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_557
timestamp 1626908933
transform 1 0 6096 0 1 333
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1073
timestamp 1626908933
transform 1 0 6720 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_503
timestamp 1626908933
transform 1 0 6720 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1042
timestamp 1626908933
transform 1 0 7776 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_412
timestamp 1626908933
transform 1 0 7776 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_501
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_242
timestamp 1626908933
transform 1 0 7488 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_611
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_243
timestamp 1626908933
transform 1 0 7584 0 -1 1332
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_104
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_374
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_104
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_374
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_104
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_374
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_111
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_399
timestamp 1626908933
transform 1 0 8600 0 1 666
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_499
timestamp 1626908933
transform 1 0 7872 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1069
timestamp 1626908933
transform 1 0 7872 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1048
timestamp 1626908933
transform 1 0 8736 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_479
timestamp 1626908933
transform 1 0 8736 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1055
timestamp 1626908933
transform 1 0 9120 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_485
timestamp 1626908933
transform 1 0 9120 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1041
timestamp 1626908933
transform 1 0 8640 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_411
timestamp 1626908933
transform 1 0 8640 0 -1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1333
timestamp 1626908933
transform 1 0 9744 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_565
timestamp 1626908933
transform 1 0 9744 0 1 555
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1028
timestamp 1626908933
transform 1 0 9888 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_459
timestamp 1626908933
transform 1 0 9888 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1042
timestamp 1626908933
transform 1 0 10464 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_472
timestamp 1626908933
transform 1 0 10464 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_610
timestamp 1626908933
transform 1 0 10272 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_242
timestamp 1626908933
transform 1 0 10272 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1003
timestamp 1626908933
transform 1 0 11328 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_434
timestamp 1626908933
transform 1 0 11328 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1040
timestamp 1626908933
transform 1 0 11232 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_410
timestamp 1626908933
transform 1 0 11232 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1021
timestamp 1626908933
transform 1 0 11712 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_451
timestamp 1626908933
transform 1 0 11712 0 -1 1332
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_95
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_383
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_359
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_89
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_359
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_89
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_359
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_89
timestamp 1626908933
transform 1 0 12600 0 1 666
box -200 -49 200 49
use L1M1_PR  L1M1_PR_631
timestamp 1626908933
transform 1 0 12816 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1419
timestamp 1626908933
transform 1 0 12816 0 1 333
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_241
timestamp 1626908933
transform 1 0 12480 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_500
timestamp 1626908933
transform 1 0 12480 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_409
timestamp 1626908933
transform 1 0 12576 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1039
timestamp 1626908933
transform 1 0 12576 0 -1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_564
timestamp 1626908933
transform 1 0 12624 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1332
timestamp 1626908933
transform 1 0 12624 0 1 555
box -32 -32 32 32
use L1M1_PR  L1M1_PR_544
timestamp 1626908933
transform 1 0 13200 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1332
timestamp 1626908933
transform 1 0 13200 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_21
timestamp 1626908933
transform 1 0 13056 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_61
timestamp 1626908933
transform 1 0 13056 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_403
timestamp 1626908933
transform 1 0 12672 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_972
timestamp 1626908933
transform 1 0 12672 0 -1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_556
timestamp 1626908933
transform 1 0 13584 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1344
timestamp 1626908933
transform 1 0 13584 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_476
timestamp 1626908933
transform 1 0 13392 0 1 555
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1244
timestamp 1626908933
transform 1 0 13392 0 1 555
box -32 -32 32 32
use L1M1_PR  L1M1_PR_543
timestamp 1626908933
transform 1 0 13392 0 1 555
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1331
timestamp 1626908933
transform 1 0 13392 0 1 555
box -29 -23 29 23
use M1M2_PR  M1M2_PR_475
timestamp 1626908933
transform 1 0 13392 0 1 999
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1243
timestamp 1626908933
transform 1 0 13392 0 1 999
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_24
timestamp 1626908933
transform 1 0 13824 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_64
timestamp 1626908933
transform 1 0 13824 0 -1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1356
timestamp 1626908933
transform 1 0 14736 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_568
timestamp 1626908933
transform 1 0 14736 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_67
timestamp 1626908933
transform 1 0 14592 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_27
timestamp 1626908933
transform 1 0 14592 0 -1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1322
timestamp 1626908933
transform 1 0 14928 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_534
timestamp 1626908933
transform 1 0 14928 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_533
timestamp 1626908933
transform 1 0 15888 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1321
timestamp 1626908933
transform 1 0 15888 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_488
timestamp 1626908933
transform 1 0 15312 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1256
timestamp 1626908933
transform 1 0 15312 0 1 333
box -32 -32 32 32
use M1M2_PR  M1M2_PR_487
timestamp 1626908933
transform 1 0 15312 0 1 777
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1255
timestamp 1626908933
transform 1 0 15312 0 1 777
box -32 -32 32 32
use L1M1_PR  L1M1_PR_555
timestamp 1626908933
transform 1 0 15312 0 1 777
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1343
timestamp 1626908933
transform 1 0 15312 0 1 777
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_30
timestamp 1626908933
transform 1 0 15360 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_70
timestamp 1626908933
transform 1 0 15360 0 -1 1332
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_74
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_344
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_74
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_344
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_74
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_344
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_367
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_79
timestamp 1626908933
transform 1 0 16600 0 1 666
box -200 -142 200 178
use L1M1_PR  L1M1_PR_528
timestamp 1626908933
transform 1 0 16560 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1316
timestamp 1626908933
transform 1 0 16560 0 1 407
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_408
timestamp 1626908933
transform 1 0 16896 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1038
timestamp 1626908933
transform 1 0 16896 0 -1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_567
timestamp 1626908933
transform 1 0 16848 0 1 999
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1355
timestamp 1626908933
transform 1 0 16848 0 1 999
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_32
timestamp 1626908933
transform 1 0 16128 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_72
timestamp 1626908933
transform 1 0 16128 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_434
timestamp 1626908933
transform 1 0 17568 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1064
timestamp 1626908933
transform 1 0 17568 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_240
timestamp 1626908933
transform 1 0 17472 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_499
timestamp 1626908933
transform 1 0 17472 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_450
timestamp 1626908933
transform 1 0 17376 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1080
timestamp 1626908933
transform 1 0 17376 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_38
timestamp 1626908933
transform 1 0 17664 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_78
timestamp 1626908933
transform 1 0 17664 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_321
timestamp 1626908933
transform 1 0 16992 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_890
timestamp 1626908933
transform 1 0 16992 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_866
timestamp 1626908933
transform 1 0 18432 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_297
timestamp 1626908933
transform 1 0 18432 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_907
timestamp 1626908933
transform 1 0 18816 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_337
timestamp 1626908933
transform 1 0 18816 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_850
timestamp 1626908933
transform 1 0 19584 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_281
timestamp 1626908933
transform 1 0 19584 0 -1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1315
timestamp 1626908933
transform 1 0 19152 0 1 407
box -29 -23 29 23
use L1M1_PR  L1M1_PR_527
timestamp 1626908933
transform 1 0 19152 0 1 407
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1392
timestamp 1626908933
transform 1 0 19056 0 1 481
box -32 -32 32 32
use M1M2_PR  M1M2_PR_624
timestamp 1626908933
transform 1 0 19056 0 1 481
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_407
timestamp 1626908933
transform 1 0 19968 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1037
timestamp 1626908933
transform 1 0 19968 0 -1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_522
timestamp 1626908933
transform 1 0 19920 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1310
timestamp 1626908933
transform 1 0 19920 0 1 333
box -29 -23 29 23
use M1M2_PR  M1M2_PR_619
timestamp 1626908933
transform 1 0 20016 0 1 925
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1387
timestamp 1626908933
transform 1 0 20016 0 1 925
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_63
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_351
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_59
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_329
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_59
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_329
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_59
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_329
timestamp 1626908933
transform 1 0 20600 0 1 666
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_309
timestamp 1626908933
transform 1 0 20064 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_879
timestamp 1626908933
transform 1 0 20064 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_830
timestamp 1626908933
transform 1 0 21024 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_261
timestamp 1626908933
transform 1 0 21024 0 -1 1332
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1306
timestamp 1626908933
transform 1 0 20976 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_518
timestamp 1626908933
transform 1 0 20976 0 1 333
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_609
timestamp 1626908933
transform 1 0 20832 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_241
timestamp 1626908933
transform 1 0 20832 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_853
timestamp 1626908933
transform 1 0 21408 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_283
timestamp 1626908933
transform 1 0 21408 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1081
timestamp 1626908933
transform 1 0 22368 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_451
timestamp 1626908933
transform 1 0 22368 0 -1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1299
timestamp 1626908933
transform 1 0 22416 0 1 333
box -29 -23 29 23
use L1M1_PR  L1M1_PR_511
timestamp 1626908933
transform 1 0 22416 0 1 333
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_627
timestamp 1626908933
transform 1 0 22176 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_259
timestamp 1626908933
transform 1 0 22176 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_833
timestamp 1626908933
transform 1 0 22656 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_263
timestamp 1626908933
transform 1 0 22656 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1036
timestamp 1626908933
transform 1 0 22560 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_406
timestamp 1626908933
transform 1 0 22560 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_498
timestamp 1626908933
transform 1 0 22464 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_239
timestamp 1626908933
transform 1 0 22464 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_798
timestamp 1626908933
transform 1 0 23424 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_229
timestamp 1626908933
transform 1 0 23424 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1035
timestamp 1626908933
transform 1 0 23808 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_405
timestamp 1626908933
transform 1 0 23808 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_810
timestamp 1626908933
transform 1 0 23904 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_240
timestamp 1626908933
transform 1 0 23904 0 -1 1332
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_335
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_47
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_314
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_44
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_314
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_44
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_314
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_44
timestamp 1626908933
transform 1 0 24600 0 1 666
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_608
timestamp 1626908933
transform 1 0 24672 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_240
timestamp 1626908933
transform 1 0 24672 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_206
timestamp 1626908933
transform 1 0 24864 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_775
timestamp 1626908933
transform 1 0 24864 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_789
timestamp 1626908933
transform 1 0 25248 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_219
timestamp 1626908933
transform 1 0 25248 0 -1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1219
timestamp 1626908933
transform 1 0 25296 0 1 407
box -32 -32 32 32
use M1M2_PR  M1M2_PR_451
timestamp 1626908933
transform 1 0 25296 0 1 407
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_761
timestamp 1626908933
transform 1 0 26016 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_192
timestamp 1626908933
transform 1 0 26016 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_767
timestamp 1626908933
transform 1 0 26496 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_197
timestamp 1626908933
transform 1 0 26496 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1034
timestamp 1626908933
transform 1 0 26400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_404
timestamp 1626908933
transform 1 0 26400 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_239
timestamp 1626908933
transform 1 0 27552 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_607
timestamp 1626908933
transform 1 0 27552 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_403
timestamp 1626908933
transform 1 0 27264 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1033
timestamp 1626908933
transform 1 0 27264 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_238
timestamp 1626908933
transform 1 0 27456 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_497
timestamp 1626908933
transform 1 0 27456 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_452
timestamp 1626908933
transform 1 0 27360 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1082
timestamp 1626908933
transform 1 0 27360 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_402
timestamp 1626908933
transform 1 0 27744 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1032
timestamp 1626908933
transform 1 0 27744 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_175
timestamp 1626908933
transform 1 0 27840 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_745
timestamp 1626908933
transform 1 0 27840 0 -1 1332
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_319
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_31
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_29
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_299
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_29
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_299
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_29
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_299
timestamp 1626908933
transform 1 0 28600 0 1 666
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_155
timestamp 1626908933
transform 1 0 28608 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_724
timestamp 1626908933
transform 1 0 28608 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1031
timestamp 1626908933
transform 1 0 28992 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_401
timestamp 1626908933
transform 1 0 28992 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_721
timestamp 1626908933
transform 1 0 29088 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_151
timestamp 1626908933
transform 1 0 29088 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1030
timestamp 1626908933
transform 1 0 29856 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_400
timestamp 1626908933
transform 1 0 29856 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_695
timestamp 1626908933
transform 1 0 29952 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_126
timestamp 1626908933
transform 1 0 29952 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_697
timestamp 1626908933
transform 1 0 30336 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_127
timestamp 1626908933
transform 1 0 30336 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_606
timestamp 1626908933
transform 1 0 31104 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_238
timestamp 1626908933
transform 1 0 31104 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_680
timestamp 1626908933
transform 1 0 31296 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_111
timestamp 1626908933
transform 1 0 31296 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_672
timestamp 1626908933
transform 1 0 31680 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_102
timestamp 1626908933
transform 1 0 31680 0 -1 1332
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_303
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_15
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_284
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_14
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_284
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_14
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_284
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_14
timestamp 1626908933
transform 1 0 32600 0 1 666
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_496
timestamp 1626908933
transform 1 0 32448 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_237
timestamp 1626908933
transform 1 0 32448 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_79
timestamp 1626908933
transform 1 0 32544 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_648
timestamp 1626908933
transform 1 0 32544 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_643
timestamp 1626908933
transform 1 0 32928 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_73
timestamp 1626908933
transform 1 0 32928 0 -1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1386
timestamp 1626908933
transform 1 0 34032 0 1 851
box -32 -32 32 32
use M1M2_PR  M1M2_PR_618
timestamp 1626908933
transform 1 0 34032 0 1 851
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1029
timestamp 1626908933
transform 1 0 33696 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_399
timestamp 1626908933
transform 1 0 33696 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_615
timestamp 1626908933
transform 1 0 33792 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_46
timestamp 1626908933
transform 1 0 33792 0 -1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_613
timestamp 1626908933
transform 1 0 34176 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_43
timestamp 1626908933
transform 1 0 34176 0 -1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_622
timestamp 1626908933
transform 1 0 35952 0 1 481
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1390
timestamp 1626908933
transform 1 0 35952 0 1 481
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_14
timestamp 1626908933
transform 1 0 34944 0 -1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_584
timestamp 1626908933
transform 1 0 34944 0 -1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1318
timestamp 1626908933
transform 1 0 144 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_530
timestamp 1626908933
transform 1 0 144 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_495
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_236
timestamp 1626908933
transform 1 0 288 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_529
timestamp 1626908933
transform 1 0 1104 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1317
timestamp 1626908933
transform 1 0 1104 0 1 1443
box -29 -23 29 23
use M1M2_PR  M1M2_PR_468
timestamp 1626908933
transform 1 0 1104 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1236
timestamp 1626908933
transform 1 0 1104 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_536
timestamp 1626908933
transform 1 0 528 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1324
timestamp 1626908933
transform 1 0 528 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_22
timestamp 1626908933
transform 1 0 1152 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_62
timestamp 1626908933
transform 1 0 1152 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_10
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_50
timestamp 1626908933
transform 1 0 384 0 1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1346
timestamp 1626908933
transform 1 0 1296 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_558
timestamp 1626908933
transform 1 0 1296 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1352
timestamp 1626908933
transform 1 0 1296 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_564
timestamp 1626908933
transform 1 0 1296 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_514
timestamp 1626908933
transform 1 0 2160 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1282
timestamp 1626908933
transform 1 0 2160 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_490
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1258
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_557
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_585
timestamp 1626908933
transform 1 0 2064 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1345
timestamp 1626908933
transform 1 0 1872 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1373
timestamp 1626908933
transform 1 0 2064 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_498
timestamp 1626908933
transform 1 0 1968 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1266
timestamp 1626908933
transform 1 0 1968 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_569
timestamp 1626908933
transform 1 0 1968 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1357
timestamp 1626908933
transform 1 0 1968 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_489
timestamp 1626908933
transform 1 0 1872 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1257
timestamp 1626908933
transform 1 0 1872 0 1 1591
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_28
timestamp 1626908933
transform 1 0 1920 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_68
timestamp 1626908933
transform 1 0 1920 0 1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_494
timestamp 1626908933
transform 1 0 2352 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1262
timestamp 1626908933
transform 1 0 2352 0 1 1073
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_269
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_539
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_269
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_539
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_269
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_539
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -49 200 49
use M1M2_PR  M1M2_PR_493
timestamp 1626908933
transform 1 0 2352 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1261
timestamp 1626908933
transform 1 0 2352 0 1 1443
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_574
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_286
timestamp 1626908933
transform 1 0 2600 0 1 1332
box -200 -142 200 178
use L1M1_PR  L1M1_PR_563
timestamp 1626908933
transform 1 0 2640 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1351
timestamp 1626908933
transform 1 0 2640 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_546
timestamp 1626908933
transform 1 0 2688 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1115
timestamp 1626908933
transform 1 0 2688 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_16
timestamp 1626908933
transform 1 0 3072 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_7
timestamp 1626908933
transform 1 0 3072 0 1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_535
timestamp 1626908933
transform 1 0 3216 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1303
timestamp 1626908933
transform 1 0 3216 0 1 1443
box -32 -32 32 32
use L1M1_PR  L1M1_PR_610
timestamp 1626908933
transform 1 0 3216 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1398
timestamp 1626908933
transform 1 0 3216 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_398
timestamp 1626908933
transform 1 0 3456 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1028
timestamp 1626908933
transform 1 0 3456 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_613
timestamp 1626908933
transform 1 0 3312 0 1 1591
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1401
timestamp 1626908933
transform 1 0 3312 0 1 1591
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_397
timestamp 1626908933
transform 1 0 3936 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1027
timestamp 1626908933
transform 1 0 3936 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_538
timestamp 1626908933
transform 1 0 3888 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1306
timestamp 1626908933
transform 1 0 3888 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_612
timestamp 1626908933
transform 1 0 3888 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1400
timestamp 1626908933
transform 1 0 3888 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_537
timestamp 1626908933
transform 1 0 3888 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1305
timestamp 1626908933
transform 1 0 3888 0 1 1591
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_533
timestamp 1626908933
transform 1 0 3552 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1102
timestamp 1626908933
transform 1 0 3552 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1113
timestamp 1626908933
transform 1 0 4032 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_543
timestamp 1626908933
transform 1 0 4032 0 1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1575
timestamp 1626908933
transform 1 0 3984 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_787
timestamp 1626908933
transform 1 0 3984 0 1 1073
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_605
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_237
timestamp 1626908933
transform 1 0 4800 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_494
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_235
timestamp 1626908933
transform 1 0 4992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_604
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_236
timestamp 1626908933
transform 1 0 5088 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1099
timestamp 1626908933
transform 1 0 5280 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_529
timestamp 1626908933
transform 1 0 5280 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_396
timestamp 1626908933
transform 1 0 6048 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1026
timestamp 1626908933
transform 1 0 6048 0 1 1332
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_558
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_270
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_524
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_254
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_524
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_254
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_524
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_254
timestamp 1626908933
transform 1 0 6600 0 1 1332
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1025
timestamp 1626908933
transform 1 0 6528 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_395
timestamp 1626908933
transform 1 0 6528 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_515
timestamp 1626908933
transform 1 0 6624 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1085
timestamp 1626908933
transform 1 0 6624 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_504
timestamp 1626908933
transform 1 0 6144 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1073
timestamp 1626908933
transform 1 0 6144 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1024
timestamp 1626908933
transform 1 0 7392 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_394
timestamp 1626908933
transform 1 0 7392 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1059
timestamp 1626908933
transform 1 0 7488 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_490
timestamp 1626908933
transform 1 0 7488 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1068
timestamp 1626908933
transform 1 0 7872 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_498
timestamp 1626908933
transform 1 0 7872 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1023
timestamp 1626908933
transform 1 0 8640 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_393
timestamp 1626908933
transform 1 0 8640 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1047
timestamp 1626908933
transform 1 0 8736 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_478
timestamp 1626908933
transform 1 0 8736 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1054
timestamp 1626908933
transform 1 0 9120 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_484
timestamp 1626908933
transform 1 0 9120 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_234
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_493
timestamp 1626908933
transform 1 0 9984 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_453
timestamp 1626908933
transform 1 0 9888 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1083
timestamp 1626908933
transform 1 0 9888 0 1 1332
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_542
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_254
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_239
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_509
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_239
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_509
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_239
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_509
timestamp 1626908933
transform 1 0 10600 0 1 1332
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_471
timestamp 1626908933
transform 1 0 10464 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1041
timestamp 1626908933
transform 1 0 10464 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_452
timestamp 1626908933
transform 1 0 10080 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1021
timestamp 1626908933
transform 1 0 10080 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1022
timestamp 1626908933
transform 1 0 11232 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_392
timestamp 1626908933
transform 1 0 11232 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1002
timestamp 1626908933
transform 1 0 11328 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_433
timestamp 1626908933
transform 1 0 11328 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1020
timestamp 1626908933
transform 1 0 11712 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_450
timestamp 1626908933
transform 1 0 11712 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_980
timestamp 1626908933
transform 1 0 12480 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_411
timestamp 1626908933
transform 1 0 12480 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1021
timestamp 1626908933
transform 1 0 12864 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_391
timestamp 1626908933
transform 1 0 12864 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1007
timestamp 1626908933
transform 1 0 12960 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_437
timestamp 1626908933
transform 1 0 12960 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_626
timestamp 1626908933
transform 1 0 13728 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1256
timestamp 1626908933
transform 1 0 13728 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1338
timestamp 1626908933
transform 1 0 13776 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_550
timestamp 1626908933
transform 1 0 13776 0 1 1221
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1250
timestamp 1626908933
transform 1 0 13968 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_482
timestamp 1626908933
transform 1 0 13968 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1387
timestamp 1626908933
transform 1 0 13968 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_599
timestamp 1626908933
transform 1 0 13968 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1357
timestamp 1626908933
transform 1 0 13872 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_589
timestamp 1626908933
transform 1 0 13872 0 1 1665
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1337
timestamp 1626908933
transform 1 0 13968 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_549
timestamp 1626908933
transform 1 0 13968 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1249
timestamp 1626908933
transform 1 0 13968 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_481
timestamp 1626908933
transform 1 0 13968 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd2_1  sky130_fd_sc_hs__dlygate4sd2_1_0
timestamp 1626908933
transform 1 0 13824 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd2_1  sky130_fd_sc_hs__dlygate4sd2_1_1
timestamp 1626908933
transform 1 0 13824 0 1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_526
timestamp 1626908933
transform 1 0 14256 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1294
timestamp 1626908933
transform 1 0 14256 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_562
timestamp 1626908933
transform 1 0 14544 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1350
timestamp 1626908933
transform 1 0 14544 0 1 1073
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_224
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_494
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_224
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_494
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_224
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_494
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_526
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_238
timestamp 1626908933
transform 1 0 14600 0 1 1332
box -200 -142 200 178
use M1M2_PR  M1M2_PR_1293
timestamp 1626908933
transform 1 0 14256 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_525
timestamp 1626908933
transform 1 0 14256 0 1 1443
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1386
timestamp 1626908933
transform 1 0 14544 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_598
timestamp 1626908933
transform 1 0 14544 0 1 1443
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_233
timestamp 1626908933
transform 1 0 14976 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_492
timestamp 1626908933
transform 1 0 14976 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_366
timestamp 1626908933
transform 1 0 14592 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_935
timestamp 1626908933
transform 1 0 14592 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_603
timestamp 1626908933
transform 1 0 15072 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_235
timestamp 1626908933
transform 1 0 15072 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_390
timestamp 1626908933
transform 1 0 15264 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1020
timestamp 1626908933
transform 1 0 15264 0 1 1332
box -38 -49 134 715
use L1M1_PR  L1M1_PR_561
timestamp 1626908933
transform 1 0 15408 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1349
timestamp 1626908933
transform 1 0 15408 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_502
timestamp 1626908933
transform 1 0 16080 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1270
timestamp 1626908933
transform 1 0 16080 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_501
timestamp 1626908933
transform 1 0 16080 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1269
timestamp 1626908933
transform 1 0 16080 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_403
timestamp 1626908933
transform 1 0 15360 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_973
timestamp 1626908933
transform 1 0 15360 0 1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_508
timestamp 1626908933
transform 1 0 16272 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1276
timestamp 1626908933
transform 1 0 16272 0 1 1073
box -32 -32 32 32
use L1M1_PR  L1M1_PR_579
timestamp 1626908933
transform 1 0 16272 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1367
timestamp 1626908933
transform 1 0 16272 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_574
timestamp 1626908933
transform 1 0 16080 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1362
timestamp 1626908933
transform 1 0 16080 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_591
timestamp 1626908933
transform 1 0 16848 0 1 1443
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1379
timestamp 1626908933
transform 1 0 16848 0 1 1443
box -29 -23 29 23
use M1M2_PR  M1M2_PR_507
timestamp 1626908933
transform 1 0 16272 0 1 1517
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1275
timestamp 1626908933
transform 1 0 16272 0 1 1517
box -32 -32 32 32
use L1M1_PR  L1M1_PR_573
timestamp 1626908933
transform 1 0 16176 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1361
timestamp 1626908933
transform 1 0 16176 0 1 1665
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_34
timestamp 1626908933
transform 1 0 16128 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_74
timestamp 1626908933
transform 1 0 16128 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_35
timestamp 1626908933
transform 1 0 16896 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_75
timestamp 1626908933
transform 1 0 16896 0 1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_590
timestamp 1626908933
transform 1 0 17712 0 1 1073
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1378
timestamp 1626908933
transform 1 0 17712 0 1 1073
box -29 -23 29 23
use M1M2_PR  M1M2_PR_518
timestamp 1626908933
transform 1 0 16944 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1286
timestamp 1626908933
transform 1 0 16944 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_517
timestamp 1626908933
transform 1 0 16944 0 1 1443
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1285
timestamp 1626908933
transform 1 0 16944 0 1 1443
box -32 -32 32 32
use L1M1_PR  L1M1_PR_578
timestamp 1626908933
transform 1 0 17616 0 1 1517
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1366
timestamp 1626908933
transform 1 0 17616 0 1 1517
box -29 -23 29 23
use L1M1_PR  L1M1_PR_583
timestamp 1626908933
transform 1 0 17040 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1371
timestamp 1626908933
transform 1 0 17040 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_512
timestamp 1626908933
transform 1 0 17424 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1280
timestamp 1626908933
transform 1 0 17424 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_37
timestamp 1626908933
transform 1 0 17664 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_77
timestamp 1626908933
transform 1 0 17664 0 1 1332
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1383
timestamp 1626908933
transform 1 0 17808 0 1 1665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_595
timestamp 1626908933
transform 1 0 17808 0 1 1665
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1290
timestamp 1626908933
transform 1 0 18288 0 1 1221
box -32 -32 32 32
use M1M2_PR  M1M2_PR_522
timestamp 1626908933
transform 1 0 18288 0 1 1221
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1382
timestamp 1626908933
transform 1 0 18384 0 1 1221
box -29 -23 29 23
use L1M1_PR  L1M1_PR_594
timestamp 1626908933
transform 1 0 18384 0 1 1221
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_222
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_510
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_479
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_209
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_479
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_209
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_479
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_209
timestamp 1626908933
transform 1 0 18600 0 1 1332
box -200 -49 200 49
use M1M2_PR  M1M2_PR_521
timestamp 1626908933
transform 1 0 18288 0 1 1665
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1289
timestamp 1626908933
transform 1 0 18288 0 1 1665
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_336
timestamp 1626908933
transform 1 0 18816 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_906
timestamp 1626908933
transform 1 0 18816 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_296
timestamp 1626908933
transform 1 0 18432 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_865
timestamp 1626908933
transform 1 0 18432 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_849
timestamp 1626908933
transform 1 0 19584 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_280
timestamp 1626908933
transform 1 0 19584 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_878
timestamp 1626908933
transform 1 0 20064 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_308
timestamp 1626908933
transform 1 0 20064 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_491
timestamp 1626908933
transform 1 0 19968 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_232
timestamp 1626908933
transform 1 0 19968 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1382
timestamp 1626908933
transform 1 0 19728 0 1 1147
box -32 -32 32 32
use M1M2_PR  M1M2_PR_614
timestamp 1626908933
transform 1 0 19728 0 1 1147
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_602
timestamp 1626908933
transform 1 0 20832 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_234
timestamp 1626908933
transform 1 0 20832 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_829
timestamp 1626908933
transform 1 0 21024 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_260
timestamp 1626908933
transform 1 0 21024 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_852
timestamp 1626908933
transform 1 0 21408 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_282
timestamp 1626908933
transform 1 0 21408 0 1 1332
box -38 -49 806 715
use M1M2_PR  M1M2_PR_587
timestamp 1626908933
transform 1 0 21744 0 1 1591
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1355
timestamp 1626908933
transform 1 0 21744 0 1 1591
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_494
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_206
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_464
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_194
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_464
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_194
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_464
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_194
timestamp 1626908933
transform 1 0 22600 0 1 1332
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1019
timestamp 1626908933
transform 1 0 22176 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_389
timestamp 1626908933
transform 1 0 22176 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_241
timestamp 1626908933
transform 1 0 22272 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_810
timestamp 1626908933
transform 1 0 22272 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_832
timestamp 1626908933
transform 1 0 22656 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_262
timestamp 1626908933
transform 1 0 22656 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_797
timestamp 1626908933
transform 1 0 23424 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_228
timestamp 1626908933
transform 1 0 23424 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1018
timestamp 1626908933
transform 1 0 23808 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_388
timestamp 1626908933
transform 1 0 23808 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_809
timestamp 1626908933
transform 1 0 23904 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_239
timestamp 1626908933
transform 1 0 23904 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_601
timestamp 1626908933
transform 1 0 25056 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_233
timestamp 1626908933
transform 1 0 25056 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_490
timestamp 1626908933
transform 1 0 24960 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_231
timestamp 1626908933
transform 1 0 24960 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_628
timestamp 1626908933
transform 1 0 24672 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_260
timestamp 1626908933
transform 1 0 24672 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1084
timestamp 1626908933
transform 1 0 24864 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_454
timestamp 1626908933
transform 1 0 24864 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_788
timestamp 1626908933
transform 1 0 25248 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_218
timestamp 1626908933
transform 1 0 25248 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_760
timestamp 1626908933
transform 1 0 26016 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_191
timestamp 1626908933
transform 1 0 26016 0 1 1332
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_478
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_190
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_449
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_179
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_449
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_179
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_449
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_179
timestamp 1626908933
transform 1 0 26600 0 1 1332
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1017
timestamp 1626908933
transform 1 0 26400 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_387
timestamp 1626908933
transform 1 0 26400 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_196
timestamp 1626908933
transform 1 0 26496 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_766
timestamp 1626908933
transform 1 0 26496 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_744
timestamp 1626908933
transform 1 0 27840 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_174
timestamp 1626908933
transform 1 0 27840 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_600
timestamp 1626908933
transform 1 0 27264 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_232
timestamp 1626908933
transform 1 0 27264 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_737
timestamp 1626908933
transform 1 0 27456 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_168
timestamp 1626908933
transform 1 0 27456 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_723
timestamp 1626908933
transform 1 0 28608 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_154
timestamp 1626908933
transform 1 0 28608 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1016
timestamp 1626908933
transform 1 0 28992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_386
timestamp 1626908933
transform 1 0 28992 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_720
timestamp 1626908933
transform 1 0 29088 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_150
timestamp 1626908933
transform 1 0 29088 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1085
timestamp 1626908933
transform 1 0 29856 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_455
timestamp 1626908933
transform 1 0 29856 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_385
timestamp 1626908933
transform 1 0 30240 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1015
timestamp 1626908933
transform 1 0 30240 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_230
timestamp 1626908933
transform 1 0 29952 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_489
timestamp 1626908933
transform 1 0 29952 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_231
timestamp 1626908933
transform 1 0 30048 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_599
timestamp 1626908933
transform 1 0 30048 0 1 1332
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_164
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_434
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_164
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_434
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_164
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_434
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_174
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_462
timestamp 1626908933
transform 1 0 30600 0 1 1332
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_126
timestamp 1626908933
transform 1 0 30336 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_696
timestamp 1626908933
transform 1 0 30336 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_598
timestamp 1626908933
transform 1 0 31104 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_230
timestamp 1626908933
transform 1 0 31104 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_679
timestamp 1626908933
transform 1 0 31296 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_110
timestamp 1626908933
transform 1 0 31296 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_671
timestamp 1626908933
transform 1 0 31680 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_101
timestamp 1626908933
transform 1 0 31680 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1014
timestamp 1626908933
transform 1 0 32448 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_384
timestamp 1626908933
transform 1 0 32448 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_647
timestamp 1626908933
transform 1 0 32544 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_78
timestamp 1626908933
transform 1 0 32544 0 1 1332
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1380
timestamp 1626908933
transform 1 0 32880 0 1 1073
box -32 -32 32 32
use M1M2_PR  M1M2_PR_612
timestamp 1626908933
transform 1 0 32880 0 1 1073
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_642
timestamp 1626908933
transform 1 0 32928 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_72
timestamp 1626908933
transform 1 0 32928 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1013
timestamp 1626908933
transform 1 0 33696 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_383
timestamp 1626908933
transform 1 0 33696 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_614
timestamp 1626908933
transform 1 0 33792 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_45
timestamp 1626908933
transform 1 0 33792 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_612
timestamp 1626908933
transform 1 0 34176 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_42
timestamp 1626908933
transform 1 0 34176 0 1 1332
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_419
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_149
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_419
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_149
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_419
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_149
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_158
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_446
timestamp 1626908933
transform 1 0 34600 0 1 1332
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_229
timestamp 1626908933
transform 1 0 34944 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_488
timestamp 1626908933
transform 1 0 34944 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_14
timestamp 1626908933
transform 1 0 35040 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_583
timestamp 1626908933
transform 1 0 35040 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_261
timestamp 1626908933
transform 1 0 35424 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_629
timestamp 1626908933
transform 1 0 35424 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_456
timestamp 1626908933
transform 1 0 35616 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1086
timestamp 1626908933
transform 1 0 35616 0 1 1332
box -38 -49 134 715
use M1M2_PR  M1M2_PR_761
timestamp 1626908933
transform 1 0 48 0 1 2183
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1529
timestamp 1626908933
transform 1 0 48 0 1 2183
box -32 -32 32 32
use L1M1_PR  L1M1_PR_783
timestamp 1626908933
transform 1 0 144 0 1 2183
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1571
timestamp 1626908933
transform 1 0 144 0 1 2183
box -29 -23 29 23
use M1M2_PR  M1M2_PR_760
timestamp 1626908933
transform 1 0 48 0 1 2479
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1528
timestamp 1626908933
transform 1 0 48 0 1 2479
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_433
timestamp 1626908933
transform 1 0 288 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1063
timestamp 1626908933
transform 1 0 288 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_759
timestamp 1626908933
transform 1 0 336 0 1 2479
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1527
timestamp 1626908933
transform 1 0 336 0 1 2479
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_430
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_142
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_403
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_133
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_403
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_133
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_403
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_133
timestamp 1626908933
transform 1 0 600 0 1 1998
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1323
timestamp 1626908933
transform 1 0 1104 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_535
timestamp 1626908933
transform 1 0 1104 0 1 2109
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1235
timestamp 1626908933
transform 1 0 1104 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_467
timestamp 1626908933
transform 1 0 1104 0 1 2109
box -32 -32 32 32
use L1M1_PR  L1M1_PR_540
timestamp 1626908933
transform 1 0 528 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1328
timestamp 1626908933
transform 1 0 528 0 1 2405
box -29 -23 29 23
use M1M2_PR  M1M2_PR_472
timestamp 1626908933
transform 1 0 1008 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1240
timestamp 1626908933
transform 1 0 1008 0 1 2405
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_19
timestamp 1626908933
transform 1 0 1152 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_59
timestamp 1626908933
transform 1 0 1152 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_13
timestamp 1626908933
transform 1 0 384 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_53
timestamp 1626908933
transform 1 0 384 0 -1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1340
timestamp 1626908933
transform 1 0 1296 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_552
timestamp 1626908933
transform 1 0 1296 0 1 2331
box -29 -23 29 23
use M1M2_PR  M1M2_PR_484
timestamp 1626908933
transform 1 0 1872 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1252
timestamp 1626908933
transform 1 0 1872 0 1 1887
box -32 -32 32 32
use L1M1_PR  L1M1_PR_551
timestamp 1626908933
transform 1 0 1872 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1339
timestamp 1626908933
transform 1 0 1872 0 1 1887
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1251
timestamp 1626908933
transform 1 0 1872 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_483
timestamp 1626908933
transform 1 0 1872 0 1 2331
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1372
timestamp 1626908933
transform 1 0 2160 0 1 2257
box -29 -23 29 23
use L1M1_PR  L1M1_PR_584
timestamp 1626908933
transform 1 0 2160 0 1 2257
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1281
timestamp 1626908933
transform 1 0 2160 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_513
timestamp 1626908933
transform 1 0 2160 0 1 2257
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1333
timestamp 1626908933
transform 1 0 1872 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_545
timestamp 1626908933
transform 1 0 1872 0 1 2553
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1246
timestamp 1626908933
transform 1 0 1872 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_478
timestamp 1626908933
transform 1 0 1872 0 1 2553
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1368
timestamp 1626908933
transform 1 0 2064 0 1 2553
box -29 -23 29 23
use L1M1_PR  L1M1_PR_580
timestamp 1626908933
transform 1 0 2064 0 1 2553
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1278
timestamp 1626908933
transform 1 0 2064 0 1 2553
box -32 -32 32 32
use M1M2_PR  M1M2_PR_510
timestamp 1626908933
transform 1 0 2064 0 1 2553
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_9
timestamp 1626908933
transform 1 0 1920 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_0
timestamp 1626908933
transform 1 0 1920 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1062
timestamp 1626908933
transform 1 0 2304 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_432
timestamp 1626908933
transform 1 0 2304 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1087
timestamp 1626908933
transform 1 0 2400 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_457
timestamp 1626908933
transform 1 0 2400 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_487
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_228
timestamp 1626908933
transform 1 0 2496 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1257
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_627
timestamp 1626908933
transform 1 0 2592 0 -1 2664
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_573
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_285
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -142 200 178
use M1M2_PR  M1M2_PR_531
timestamp 1626908933
transform 1 0 2928 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1299
timestamp 1626908933
transform 1 0 2928 0 1 2109
box -32 -32 32 32
use L1M1_PR  L1M1_PR_606
timestamp 1626908933
transform 1 0 2832 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1394
timestamp 1626908933
transform 1 0 2832 0 1 2109
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_5
timestamp 1626908933
transform 1 0 2688 0 -1 2664
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_2
timestamp 1626908933
transform 1 0 2688 0 -1 2664
box -38 -49 614 715
use L1M1_PR  L1M1_PR_1396
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -29 -23 29 23
use L1M1_PR  L1M1_PR_608
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1301
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -32 -32 32 32
use M1M2_PR  M1M2_PR_533
timestamp 1626908933
transform 1 0 3120 0 1 2405
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1115
timestamp 1626908933
transform 1 0 3360 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_545
timestamp 1626908933
transform 1 0 3360 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1258
timestamp 1626908933
transform 1 0 3264 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_628
timestamp 1626908933
transform 1 0 3264 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1012
timestamp 1626908933
transform 1 0 4128 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_382
timestamp 1626908933
transform 1 0 4128 0 -1 2664
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_118
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_388
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_118
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_388
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_118
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_388
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_126
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_414
timestamp 1626908933
transform 1 0 4600 0 1 1998
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_532
timestamp 1626908933
transform 1 0 4608 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1102
timestamp 1626908933
transform 1 0 4608 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_522
timestamp 1626908933
transform 1 0 4224 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1091
timestamp 1626908933
transform 1 0 4224 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_597
timestamp 1626908933
transform 1 0 5760 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_229
timestamp 1626908933
transform 1 0 5760 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1085
timestamp 1626908933
transform 1 0 5376 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_516
timestamp 1626908933
transform 1 0 5376 0 -1 2664
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_557
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_269
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1087
timestamp 1626908933
transform 1 0 5952 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_517
timestamp 1626908933
transform 1 0 5952 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1072
timestamp 1626908933
transform 1 0 6720 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_502
timestamp 1626908933
transform 1 0 6720 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1011
timestamp 1626908933
transform 1 0 7776 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_381
timestamp 1626908933
transform 1 0 7776 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_596
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_228
timestamp 1626908933
transform 1 0 7584 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_486
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_227
timestamp 1626908933
transform 1 0 7488 0 -1 2664
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_103
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_373
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_103
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_373
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_103
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_373
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_110
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_398
timestamp 1626908933
transform 1 0 8600 0 1 1998
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_497
timestamp 1626908933
transform 1 0 7872 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1067
timestamp 1626908933
transform 1 0 7872 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1046
timestamp 1626908933
transform 1 0 8736 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_477
timestamp 1626908933
transform 1 0 8736 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1053
timestamp 1626908933
transform 1 0 9120 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_483
timestamp 1626908933
transform 1 0 9120 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1010
timestamp 1626908933
transform 1 0 8640 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_380
timestamp 1626908933
transform 1 0 8640 0 -1 2664
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_253
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_541
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1027
timestamp 1626908933
transform 1 0 9888 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_458
timestamp 1626908933
transform 1 0 9888 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_595
timestamp 1626908933
transform 1 0 10272 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_227
timestamp 1626908933
transform 1 0 10272 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1040
timestamp 1626908933
transform 1 0 10464 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_470
timestamp 1626908933
transform 1 0 10464 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1009
timestamp 1626908933
transform 1 0 11232 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_379
timestamp 1626908933
transform 1 0 11232 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1001
timestamp 1626908933
transform 1 0 11328 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_432
timestamp 1626908933
transform 1 0 11328 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1019
timestamp 1626908933
transform 1 0 11712 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_449
timestamp 1626908933
transform 1 0 11712 0 -1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_382
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_94
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_358
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_88
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_358
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_88
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_358
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_88
timestamp 1626908933
transform 1 0 12600 0 1 1998
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_971
timestamp 1626908933
transform 1 0 12576 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_402
timestamp 1626908933
transform 1 0 12576 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_485
timestamp 1626908933
transform 1 0 12480 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_226
timestamp 1626908933
transform 1 0 12480 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1006
timestamp 1626908933
transform 1 0 12960 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_436
timestamp 1626908933
transform 1 0 12960 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_953
timestamp 1626908933
transform 1 0 13920 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_384
timestamp 1626908933
transform 1 0 13920 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_594
timestamp 1626908933
transform 1 0 13728 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_226
timestamp 1626908933
transform 1 0 13728 0 -1 2664
box -38 -49 230 715
use osc_core_VIA4  osc_core_VIA4_237
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_525
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_992
timestamp 1626908933
transform 1 0 14304 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_422
timestamp 1626908933
transform 1 0 14304 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1008
timestamp 1626908933
transform 1 0 15072 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_378
timestamp 1626908933
transform 1 0 15072 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_934
timestamp 1626908933
transform 1 0 15168 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_365
timestamp 1626908933
transform 1 0 15168 0 -1 2664
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1360
timestamp 1626908933
transform 1 0 15504 0 1 2257
box -32 -32 32 32
use M1M2_PR  M1M2_PR_592
timestamp 1626908933
transform 1 0 15504 0 1 2257
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_972
timestamp 1626908933
transform 1 0 15552 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_402
timestamp 1626908933
transform 1 0 15552 0 -1 2664
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_73
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_343
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_73
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_343
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_73
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_343
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_78
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_366
timestamp 1626908933
transform 1 0 16600 0 1 1998
box -200 -142 200 178
use L1M1_PR  L1M1_PR_587
timestamp 1626908933
transform 1 0 16848 0 1 2331
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1375
timestamp 1626908933
transform 1 0 16848 0 1 2331
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_340
timestamp 1626908933
transform 1 0 16320 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_909
timestamp 1626908933
transform 1 0 16320 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_36
timestamp 1626908933
transform 1 0 16704 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_76
timestamp 1626908933
transform 1 0 16704 0 -1 2664
box -38 -49 806 715
use M1M2_PR  M1M2_PR_516
timestamp 1626908933
transform 1 0 16944 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1284
timestamp 1626908933
transform 1 0 16944 0 1 1887
box -32 -32 32 32
use M1M2_PR  M1M2_PR_515
timestamp 1626908933
transform 1 0 16944 0 1 2331
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1283
timestamp 1626908933
transform 1 0 16944 0 1 2331
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_225
timestamp 1626908933
transform 1 0 17568 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_593
timestamp 1626908933
transform 1 0 17568 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_225
timestamp 1626908933
transform 1 0 17472 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_484
timestamp 1626908933
transform 1 0 17472 0 -1 2664
box -38 -49 134 715
use M1M2_PR  M1M2_PR_511
timestamp 1626908933
transform 1 0 17424 0 1 2109
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1279
timestamp 1626908933
transform 1 0 17424 0 1 2109
box -32 -32 32 32
use L1M1_PR  L1M1_PR_582
timestamp 1626908933
transform 1 0 17424 0 1 2109
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1370
timestamp 1626908933
transform 1 0 17424 0 1 2109
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_315
timestamp 1626908933
transform 1 0 17760 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_884
timestamp 1626908933
transform 1 0 17760 0 -1 2664
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_221
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_509
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_923
timestamp 1626908933
transform 1 0 18144 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_353
timestamp 1626908933
transform 1 0 18144 0 -1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1374
timestamp 1626908933
transform 1 0 18384 0 1 1887
box -29 -23 29 23
use L1M1_PR  L1M1_PR_586
timestamp 1626908933
transform 1 0 18384 0 1 1887
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_860
timestamp 1626908933
transform 1 0 18912 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_291
timestamp 1626908933
transform 1 0 18912 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1007
timestamp 1626908933
transform 1 0 19296 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_377
timestamp 1626908933
transform 1 0 19296 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_901
timestamp 1626908933
transform 1 0 19392 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_331
timestamp 1626908933
transform 1 0 19392 0 -1 2664
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_328
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_58
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_328
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_58
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_328
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_58
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_62
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_350
timestamp 1626908933
transform 1 0 20600 0 1 1998
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_592
timestamp 1626908933
transform 1 0 20160 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_224
timestamp 1626908933
transform 1 0 20160 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_275
timestamp 1626908933
transform 1 0 20352 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_844
timestamp 1626908933
transform 1 0 20352 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_866
timestamp 1626908933
transform 1 0 20736 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_296
timestamp 1626908933
transform 1 0 20736 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_591
timestamp 1626908933
transform 1 0 21504 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_223
timestamp 1626908933
transform 1 0 21504 0 -1 2664
box -38 -49 230 715
use osc_core_VIA4  osc_core_VIA4_493
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_205
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -142 200 178
use M1M2_PR  M1M2_PR_1358
timestamp 1626908933
transform 1 0 22320 0 1 2183
box -32 -32 32 32
use M1M2_PR  M1M2_PR_590
timestamp 1626908933
transform 1 0 22320 0 1 2183
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_842
timestamp 1626908933
transform 1 0 21696 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_272
timestamp 1626908933
transform 1 0 21696 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1006
timestamp 1626908933
transform 1 0 22560 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_376
timestamp 1626908933
transform 1 0 22560 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_831
timestamp 1626908933
transform 1 0 22656 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_261
timestamp 1626908933
transform 1 0 22656 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_483
timestamp 1626908933
transform 1 0 22464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_224
timestamp 1626908933
transform 1 0 22464 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_796
timestamp 1626908933
transform 1 0 23424 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_227
timestamp 1626908933
transform 1 0 23424 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1005
timestamp 1626908933
transform 1 0 23808 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_375
timestamp 1626908933
transform 1 0 23808 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_808
timestamp 1626908933
transform 1 0 23904 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_238
timestamp 1626908933
transform 1 0 23904 0 -1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_334
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_46
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_313
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_43
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_313
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_43
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_313
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_43
timestamp 1626908933
transform 1 0 24600 0 1 1998
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_590
timestamp 1626908933
transform 1 0 24672 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_222
timestamp 1626908933
transform 1 0 24672 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_205
timestamp 1626908933
transform 1 0 24864 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_774
timestamp 1626908933
transform 1 0 24864 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_787
timestamp 1626908933
transform 1 0 25248 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_217
timestamp 1626908933
transform 1 0 25248 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_759
timestamp 1626908933
transform 1 0 26016 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_190
timestamp 1626908933
transform 1 0 26016 0 -1 2664
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_477
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_189
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1004
timestamp 1626908933
transform 1 0 26400 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_374
timestamp 1626908933
transform 1 0 26400 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_765
timestamp 1626908933
transform 1 0 26496 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_195
timestamp 1626908933
transform 1 0 26496 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_221
timestamp 1626908933
transform 1 0 27552 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_589
timestamp 1626908933
transform 1 0 27552 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_223
timestamp 1626908933
transform 1 0 27456 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_482
timestamp 1626908933
transform 1 0 27456 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_373
timestamp 1626908933
transform 1 0 27264 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_458
timestamp 1626908933
transform 1 0 27360 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1003
timestamp 1626908933
transform 1 0 27264 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1088
timestamp 1626908933
transform 1 0 27360 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_372
timestamp 1626908933
transform 1 0 27744 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1002
timestamp 1626908933
transform 1 0 27744 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_173
timestamp 1626908933
transform 1 0 27840 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_743
timestamp 1626908933
transform 1 0 27840 0 -1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_318
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_30
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_28
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_298
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_28
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_298
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_28
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_298
timestamp 1626908933
transform 1 0 28600 0 1 1998
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_153
timestamp 1626908933
transform 1 0 28608 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_722
timestamp 1626908933
transform 1 0 28608 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1001
timestamp 1626908933
transform 1 0 28992 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_371
timestamp 1626908933
transform 1 0 28992 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_719
timestamp 1626908933
transform 1 0 29088 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_149
timestamp 1626908933
transform 1 0 29088 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1000
timestamp 1626908933
transform 1 0 29856 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_370
timestamp 1626908933
transform 1 0 29856 0 -1 2664
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_461
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_173
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_694
timestamp 1626908933
transform 1 0 29952 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_125
timestamp 1626908933
transform 1 0 29952 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_695
timestamp 1626908933
transform 1 0 30336 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_125
timestamp 1626908933
transform 1 0 30336 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_588
timestamp 1626908933
transform 1 0 31104 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_220
timestamp 1626908933
transform 1 0 31104 0 -1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_678
timestamp 1626908933
transform 1 0 31296 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_109
timestamp 1626908933
transform 1 0 31296 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_670
timestamp 1626908933
transform 1 0 31680 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_100
timestamp 1626908933
transform 1 0 31680 0 -1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_302
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_14
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_283
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_13
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_283
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_13
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_283
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_13
timestamp 1626908933
transform 1 0 32600 0 1 1998
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_481
timestamp 1626908933
transform 1 0 32448 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_222
timestamp 1626908933
transform 1 0 32448 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_77
timestamp 1626908933
transform 1 0 32544 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_646
timestamp 1626908933
transform 1 0 32544 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_641
timestamp 1626908933
transform 1 0 32928 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_71
timestamp 1626908933
transform 1 0 32928 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_999
timestamp 1626908933
transform 1 0 33696 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_369
timestamp 1626908933
transform 1 0 33696 0 -1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_613
timestamp 1626908933
transform 1 0 33792 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_44
timestamp 1626908933
transform 1 0 33792 0 -1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_611
timestamp 1626908933
transform 1 0 34176 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_41
timestamp 1626908933
transform 1 0 34176 0 -1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_157
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_445
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_13
timestamp 1626908933
transform 1 0 34944 0 -1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_583
timestamp 1626908933
transform 1 0 34944 0 -1 2664
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1334
timestamp 1626908933
transform 1 0 528 0 1 2923
box -29 -23 29 23
use L1M1_PR  L1M1_PR_546
timestamp 1626908933
transform 1 0 528 0 1 2923
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_429
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_141
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_402
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_132
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_402
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_132
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_402
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_132
timestamp 1626908933
transform 1 0 600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_979
timestamp 1626908933
transform 1 0 288 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_349
timestamp 1626908933
transform 1 0 288 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_480
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_221
timestamp 1626908933
transform 1 0 288 0 1 2664
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1327
timestamp 1626908933
transform 1 0 1104 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_539
timestamp 1626908933
transform 1 0 1104 0 1 2775
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1239
timestamp 1626908933
transform 1 0 1008 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_471
timestamp 1626908933
transform 1 0 1008 0 1 2775
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1364
timestamp 1626908933
transform 1 0 1200 0 1 2997
box -29 -23 29 23
use L1M1_PR  L1M1_PR_576
timestamp 1626908933
transform 1 0 1200 0 1 2997
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1272
timestamp 1626908933
transform 1 0 1296 0 1 2997
box -32 -32 32 32
use M1M2_PR  M1M2_PR_504
timestamp 1626908933
transform 1 0 1296 0 1 2997
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_1
timestamp 1626908933
transform 1 0 1152 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_4
timestamp 1626908933
transform 1 0 1152 0 -1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_16
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_56
timestamp 1626908933
transform 1 0 384 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_569
timestamp 1626908933
transform 1 0 384 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1139
timestamp 1626908933
transform 1 0 384 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__bufbuf_8  sky130_fd_sc_hs__bufbuf_8_1
timestamp 1626908933
transform 1 0 1152 0 1 2664
box -38 -49 1478 715
use sky130_fd_sc_hs__bufbuf_8  sky130_fd_sc_hs__bufbuf_8_0
timestamp 1626908933
transform 1 0 1152 0 1 2664
box -38 -49 1478 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1127
timestamp 1626908933
transform 1 0 1728 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_557
timestamp 1626908933
transform 1 0 1728 0 -1 3996
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1358
timestamp 1626908933
transform 1 0 1872 0 1 2775
box -29 -23 29 23
use L1M1_PR  L1M1_PR_570
timestamp 1626908933
transform 1 0 1872 0 1 2775
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1265
timestamp 1626908933
transform 1 0 1968 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_497
timestamp 1626908933
transform 1 0 1968 0 1 2775
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1245
timestamp 1626908933
transform 1 0 1872 0 1 2923
box -32 -32 32 32
use M1M2_PR  M1M2_PR_477
timestamp 1626908933
transform 1 0 1872 0 1 2923
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_538
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_268
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_538
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_268
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_538
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_268
timestamp 1626908933
transform 1 0 2600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_472
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_213
timestamp 1626908933
transform 1 0 2496 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_978
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_348
timestamp 1626908933
transform 1 0 2592 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1259
timestamp 1626908933
transform 1 0 2592 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_629
timestamp 1626908933
transform 1 0 2592 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_551
timestamp 1626908933
transform 1 0 2688 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1121
timestamp 1626908933
transform 1 0 2688 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_550
timestamp 1626908933
transform 1 0 2688 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1120
timestamp 1626908933
transform 1 0 2688 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_368
timestamp 1626908933
transform 1 0 3456 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_998
timestamp 1626908933
transform 1 0 3456 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_347
timestamp 1626908933
transform 1 0 3456 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_977
timestamp 1626908933
transform 1 0 3456 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_367
timestamp 1626908933
transform 1 0 3936 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_997
timestamp 1626908933
transform 1 0 3936 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_346
timestamp 1626908933
transform 1 0 3936 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_976
timestamp 1626908933
transform 1 0 3936 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_532
timestamp 1626908933
transform 1 0 3552 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1101
timestamp 1626908933
transform 1 0 3552 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_531
timestamp 1626908933
transform 1 0 3552 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1100
timestamp 1626908933
transform 1 0 3552 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1111
timestamp 1626908933
transform 1 0 4032 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_541
timestamp 1626908933
transform 1 0 4032 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1112
timestamp 1626908933
transform 1 0 4032 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_542
timestamp 1626908933
transform 1 0 4032 0 1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_413
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_125
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_117
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_387
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_117
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_387
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_117
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_387
timestamp 1626908933
transform 1 0 4600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_220
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_479
timestamp 1626908933
transform 1 0 4992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_219
timestamp 1626908933
transform 1 0 4800 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_587
timestamp 1626908933
transform 1 0 4800 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_345
timestamp 1626908933
transform 1 0 4800 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_975
timestamp 1626908933
transform 1 0 4800 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_520
timestamp 1626908933
transform 1 0 4896 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1089
timestamp 1626908933
transform 1 0 4896 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1097
timestamp 1626908933
transform 1 0 5280 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_527
timestamp 1626908933
transform 1 0 5280 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_586
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_218
timestamp 1626908933
transform 1 0 5088 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1098
timestamp 1626908933
transform 1 0 5280 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_528
timestamp 1626908933
transform 1 0 5280 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_366
timestamp 1626908933
transform 1 0 6048 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_996
timestamp 1626908933
transform 1 0 6048 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_344
timestamp 1626908933
transform 1 0 6048 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_974
timestamp 1626908933
transform 1 0 6048 0 -1 3996
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_523
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_253
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_523
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_253
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_523
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_253
timestamp 1626908933
transform 1 0 6600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_973
timestamp 1626908933
transform 1 0 6528 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_343
timestamp 1626908933
transform 1 0 6528 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_995
timestamp 1626908933
transform 1 0 6528 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_365
timestamp 1626908933
transform 1 0 6528 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_514
timestamp 1626908933
transform 1 0 6624 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1084
timestamp 1626908933
transform 1 0 6624 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_503
timestamp 1626908933
transform 1 0 6144 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1072
timestamp 1626908933
transform 1 0 6144 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_513
timestamp 1626908933
transform 1 0 6624 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1083
timestamp 1626908933
transform 1 0 6624 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_502
timestamp 1626908933
transform 1 0 6144 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1071
timestamp 1626908933
transform 1 0 6144 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1093
timestamp 1626908933
transform 1 0 7392 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_463
timestamp 1626908933
transform 1 0 7392 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_471
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_212
timestamp 1626908933
transform 1 0 7488 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_994
timestamp 1626908933
transform 1 0 7392 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_364
timestamp 1626908933
transform 1 0 7392 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_972
timestamp 1626908933
transform 1 0 7776 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_342
timestamp 1626908933
transform 1 0 7776 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_578
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_210
timestamp 1626908933
transform 1 0 7584 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_489
timestamp 1626908933
transform 1 0 7488 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1058
timestamp 1626908933
transform 1 0 7488 0 1 2664
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_102
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_372
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_102
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_372
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_102
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_372
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_109
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_397
timestamp 1626908933
transform 1 0 8600 0 1 3330
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_496
timestamp 1626908933
transform 1 0 7872 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1066
timestamp 1626908933
transform 1 0 7872 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_495
timestamp 1626908933
transform 1 0 7872 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1065
timestamp 1626908933
transform 1 0 7872 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_363
timestamp 1626908933
transform 1 0 8640 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_993
timestamp 1626908933
transform 1 0 8640 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_341
timestamp 1626908933
transform 1 0 8640 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_971
timestamp 1626908933
transform 1 0 8640 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_482
timestamp 1626908933
transform 1 0 9120 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1052
timestamp 1626908933
transform 1 0 9120 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_476
timestamp 1626908933
transform 1 0 8736 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1045
timestamp 1626908933
transform 1 0 8736 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_481
timestamp 1626908933
transform 1 0 9120 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1051
timestamp 1626908933
transform 1 0 9120 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_475
timestamp 1626908933
transform 1 0 8736 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1044
timestamp 1626908933
transform 1 0 8736 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_219
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_478
timestamp 1626908933
transform 1 0 9984 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_459
timestamp 1626908933
transform 1 0 9888 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1089
timestamp 1626908933
transform 1 0 9888 0 1 2664
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_238
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_508
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_238
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_508
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_238
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_508
timestamp 1626908933
transform 1 0 10600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_209
timestamp 1626908933
transform 1 0 10272 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_577
timestamp 1626908933
transform 1 0 10272 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_469
timestamp 1626908933
transform 1 0 10464 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1039
timestamp 1626908933
transform 1 0 10464 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_451
timestamp 1626908933
transform 1 0 10080 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1020
timestamp 1626908933
transform 1 0 10080 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_468
timestamp 1626908933
transform 1 0 10464 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1038
timestamp 1626908933
transform 1 0 10464 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_457
timestamp 1626908933
transform 1 0 9888 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1026
timestamp 1626908933
transform 1 0 9888 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_970
timestamp 1626908933
transform 1 0 11232 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_340
timestamp 1626908933
transform 1 0 11232 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_999
timestamp 1626908933
transform 1 0 11328 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_430
timestamp 1626908933
transform 1 0 11328 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_992
timestamp 1626908933
transform 1 0 11232 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_362
timestamp 1626908933
transform 1 0 11232 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1000
timestamp 1626908933
transform 1 0 11328 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_431
timestamp 1626908933
transform 1 0 11328 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1017
timestamp 1626908933
transform 1 0 11712 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_447
timestamp 1626908933
transform 1 0 11712 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1018
timestamp 1626908933
transform 1 0 11712 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_448
timestamp 1626908933
transform 1 0 11712 0 1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_381
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_93
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_357
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_87
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_357
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_87
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_357
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_87
timestamp 1626908933
transform 1 0 12600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_361
timestamp 1626908933
transform 1 0 12864 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_991
timestamp 1626908933
transform 1 0 12864 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_211
timestamp 1626908933
transform 1 0 12480 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_470
timestamp 1626908933
transform 1 0 12480 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_435
timestamp 1626908933
transform 1 0 12960 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1005
timestamp 1626908933
transform 1 0 12960 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_410
timestamp 1626908933
transform 1 0 12480 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_979
timestamp 1626908933
transform 1 0 12480 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_434
timestamp 1626908933
transform 1 0 12960 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1004
timestamp 1626908933
transform 1 0 12960 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_401
timestamp 1626908933
transform 1 0 12576 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_970
timestamp 1626908933
transform 1 0 12576 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_951
timestamp 1626908933
transform 1 0 13920 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_382
timestamp 1626908933
transform 1 0 13920 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_576
timestamp 1626908933
transform 1 0 13728 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_208
timestamp 1626908933
transform 1 0 13728 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_990
timestamp 1626908933
transform 1 0 13728 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_360
timestamp 1626908933
transform 1 0 13728 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_952
timestamp 1626908933
transform 1 0 13824 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_383
timestamp 1626908933
transform 1 0 13824 0 1 2664
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_223
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_493
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_223
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_493
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_223
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_493
timestamp 1626908933
transform 1 0 14600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_218
timestamp 1626908933
transform 1 0 14976 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_477
timestamp 1626908933
transform 1 0 14976 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_421
timestamp 1626908933
transform 1 0 14208 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_991
timestamp 1626908933
transform 1 0 14208 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_420
timestamp 1626908933
transform 1 0 14304 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_990
timestamp 1626908933
transform 1 0 14304 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_969
timestamp 1626908933
transform 1 0 15072 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_339
timestamp 1626908933
transform 1 0 15072 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_932
timestamp 1626908933
transform 1 0 15168 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_363
timestamp 1626908933
transform 1 0 15168 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_989
timestamp 1626908933
transform 1 0 15072 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_359
timestamp 1626908933
transform 1 0 15072 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_933
timestamp 1626908933
transform 1 0 15168 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_364
timestamp 1626908933
transform 1 0 15168 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_970
timestamp 1626908933
transform 1 0 15552 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_400
timestamp 1626908933
transform 1 0 15552 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_971
timestamp 1626908933
transform 1 0 15552 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_401
timestamp 1626908933
transform 1 0 15552 0 1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_365
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_77
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_342
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_72
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_342
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_72
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_342
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_72
timestamp 1626908933
transform 1 0 16600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_585
timestamp 1626908933
transform 1 0 16320 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_217
timestamp 1626908933
transform 1 0 16320 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_339
timestamp 1626908933
transform 1 0 16512 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_908
timestamp 1626908933
transform 1 0 16512 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_375
timestamp 1626908933
transform 1 0 16896 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_945
timestamp 1626908933
transform 1 0 16896 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_338
timestamp 1626908933
transform 1 0 16320 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_907
timestamp 1626908933
transform 1 0 16320 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_374
timestamp 1626908933
transform 1 0 16704 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_944
timestamp 1626908933
transform 1 0 16704 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_358
timestamp 1626908933
transform 1 0 17664 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_988
timestamp 1626908933
transform 1 0 17664 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_207
timestamp 1626908933
transform 1 0 17568 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_575
timestamp 1626908933
transform 1 0 17568 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_210
timestamp 1626908933
transform 1 0 17472 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_469
timestamp 1626908933
transform 1 0 17472 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_314
timestamp 1626908933
transform 1 0 17760 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_883
timestamp 1626908933
transform 1 0 17760 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_313
timestamp 1626908933
transform 1 0 17760 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_882
timestamp 1626908933
transform 1 0 17760 0 -1 3996
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_208
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_478
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_208
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_478
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_208
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_478
timestamp 1626908933
transform 1 0 18600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_352
timestamp 1626908933
transform 1 0 18144 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_922
timestamp 1626908933
transform 1 0 18144 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_351
timestamp 1626908933
transform 1 0 18144 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_921
timestamp 1626908933
transform 1 0 18144 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_216
timestamp 1626908933
transform 1 0 18912 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_584
timestamp 1626908933
transform 1 0 18912 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_357
timestamp 1626908933
transform 1 0 19104 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_987
timestamp 1626908933
transform 1 0 19104 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_338
timestamp 1626908933
transform 1 0 19296 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_968
timestamp 1626908933
transform 1 0 19296 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_330
timestamp 1626908933
transform 1 0 19200 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_900
timestamp 1626908933
transform 1 0 19200 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_329
timestamp 1626908933
transform 1 0 19392 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_899
timestamp 1626908933
transform 1 0 19392 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_290
timestamp 1626908933
transform 1 0 18912 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_859
timestamp 1626908933
transform 1 0 18912 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_217
timestamp 1626908933
transform 1 0 19968 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_476
timestamp 1626908933
transform 1 0 19968 0 1 2664
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_327
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_57
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_327
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_57
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_327
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_57
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_61
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_349
timestamp 1626908933
transform 1 0 20600 0 1 3330
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_574
timestamp 1626908933
transform 1 0 20160 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_206
timestamp 1626908933
transform 1 0 20160 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_307
timestamp 1626908933
transform 1 0 20064 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_877
timestamp 1626908933
transform 1 0 20064 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_274
timestamp 1626908933
transform 1 0 20352 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_843
timestamp 1626908933
transform 1 0 20352 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_865
timestamp 1626908933
transform 1 0 20736 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_295
timestamp 1626908933
transform 1 0 20736 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_573
timestamp 1626908933
transform 1 0 21504 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_205
timestamp 1626908933
transform 1 0 21504 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_583
timestamp 1626908933
transform 1 0 20832 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_215
timestamp 1626908933
transform 1 0 20832 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_828
timestamp 1626908933
transform 1 0 21024 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_259
timestamp 1626908933
transform 1 0 21024 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_851
timestamp 1626908933
transform 1 0 21408 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_281
timestamp 1626908933
transform 1 0 21408 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_356
timestamp 1626908933
transform 1 0 22176 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_986
timestamp 1626908933
transform 1 0 22176 0 1 2664
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_193
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_463
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_193
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_463
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_193
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_463
timestamp 1626908933
transform 1 0 22600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_240
timestamp 1626908933
transform 1 0 22272 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_809
timestamp 1626908933
transform 1 0 22272 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_271
timestamp 1626908933
transform 1 0 21696 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_841
timestamp 1626908933
transform 1 0 21696 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_967
timestamp 1626908933
transform 1 0 22560 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_337
timestamp 1626908933
transform 1 0 22560 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_829
timestamp 1626908933
transform 1 0 22656 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_259
timestamp 1626908933
transform 1 0 22656 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_468
timestamp 1626908933
transform 1 0 22464 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_209
timestamp 1626908933
transform 1 0 22464 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_830
timestamp 1626908933
transform 1 0 22656 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_260
timestamp 1626908933
transform 1 0 22656 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_794
timestamp 1626908933
transform 1 0 23424 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_225
timestamp 1626908933
transform 1 0 23424 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_795
timestamp 1626908933
transform 1 0 23424 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_226
timestamp 1626908933
transform 1 0 23424 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_966
timestamp 1626908933
transform 1 0 23808 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_336
timestamp 1626908933
transform 1 0 23808 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_806
timestamp 1626908933
transform 1 0 23904 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_236
timestamp 1626908933
transform 1 0 23904 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_985
timestamp 1626908933
transform 1 0 23808 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_355
timestamp 1626908933
transform 1 0 23808 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_807
timestamp 1626908933
transform 1 0 23904 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_237
timestamp 1626908933
transform 1 0 23904 0 1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_333
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_45
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_312
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_42
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_312
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_42
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_312
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_42
timestamp 1626908933
transform 1 0 24600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_572
timestamp 1626908933
transform 1 0 24672 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_204
timestamp 1626908933
transform 1 0 24672 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_630
timestamp 1626908933
transform 1 0 24672 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_262
timestamp 1626908933
transform 1 0 24672 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_460
timestamp 1626908933
transform 1 0 24864 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1090
timestamp 1626908933
transform 1 0 24864 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_216
timestamp 1626908933
transform 1 0 24960 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_475
timestamp 1626908933
transform 1 0 24960 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_214
timestamp 1626908933
transform 1 0 25056 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_582
timestamp 1626908933
transform 1 0 25056 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_204
timestamp 1626908933
transform 1 0 24864 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_773
timestamp 1626908933
transform 1 0 24864 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_785
timestamp 1626908933
transform 1 0 25248 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_215
timestamp 1626908933
transform 1 0 25248 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_757
timestamp 1626908933
transform 1 0 26016 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_188
timestamp 1626908933
transform 1 0 26016 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_786
timestamp 1626908933
transform 1 0 25248 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_216
timestamp 1626908933
transform 1 0 25248 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_758
timestamp 1626908933
transform 1 0 26016 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_189
timestamp 1626908933
transform 1 0 26016 0 1 2664
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_448
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_178
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_448
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_178
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_448
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_178
timestamp 1626908933
transform 1 0 26600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_965
timestamp 1626908933
transform 1 0 26400 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_335
timestamp 1626908933
transform 1 0 26400 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_984
timestamp 1626908933
transform 1 0 26400 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_354
timestamp 1626908933
transform 1 0 26400 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_194
timestamp 1626908933
transform 1 0 26496 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_764
timestamp 1626908933
transform 1 0 26496 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_193
timestamp 1626908933
transform 1 0 26496 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_763
timestamp 1626908933
transform 1 0 26496 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_964
timestamp 1626908933
transform 1 0 27264 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_334
timestamp 1626908933
transform 1 0 27264 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1094
timestamp 1626908933
transform 1 0 27360 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_464
timestamp 1626908933
transform 1 0 27360 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_467
timestamp 1626908933
transform 1 0 27456 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_208
timestamp 1626908933
transform 1 0 27456 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_571
timestamp 1626908933
transform 1 0 27552 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_203
timestamp 1626908933
transform 1 0 27552 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_581
timestamp 1626908933
transform 1 0 27264 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_213
timestamp 1626908933
transform 1 0 27264 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_333
timestamp 1626908933
transform 1 0 27744 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_963
timestamp 1626908933
transform 1 0 27744 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_167
timestamp 1626908933
transform 1 0 27456 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_736
timestamp 1626908933
transform 1 0 27456 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_172
timestamp 1626908933
transform 1 0 27840 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_742
timestamp 1626908933
transform 1 0 27840 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_171
timestamp 1626908933
transform 1 0 27840 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_741
timestamp 1626908933
transform 1 0 27840 0 -1 3996
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_317
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_29
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_27
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_297
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_27
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_297
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_27
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_297
timestamp 1626908933
transform 1 0 28600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_152
timestamp 1626908933
transform 1 0 28608 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_721
timestamp 1626908933
transform 1 0 28608 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_151
timestamp 1626908933
transform 1 0 28608 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_720
timestamp 1626908933
transform 1 0 28608 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_962
timestamp 1626908933
transform 1 0 28992 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_332
timestamp 1626908933
transform 1 0 28992 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_983
timestamp 1626908933
transform 1 0 28992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_353
timestamp 1626908933
transform 1 0 28992 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_717
timestamp 1626908933
transform 1 0 29088 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_147
timestamp 1626908933
transform 1 0 29088 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_961
timestamp 1626908933
transform 1 0 29856 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_331
timestamp 1626908933
transform 1 0 29856 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_718
timestamp 1626908933
transform 1 0 29088 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_148
timestamp 1626908933
transform 1 0 29088 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1091
timestamp 1626908933
transform 1 0 29856 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_461
timestamp 1626908933
transform 1 0 29856 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_352
timestamp 1626908933
transform 1 0 30240 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_982
timestamp 1626908933
transform 1 0 30240 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_215
timestamp 1626908933
transform 1 0 29952 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_474
timestamp 1626908933
transform 1 0 29952 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_212
timestamp 1626908933
transform 1 0 30048 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_580
timestamp 1626908933
transform 1 0 30048 0 1 2664
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_163
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_433
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_163
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_433
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_163
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_433
timestamp 1626908933
transform 1 0 30600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_124
timestamp 1626908933
transform 1 0 30336 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_694
timestamp 1626908933
transform 1 0 30336 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_123
timestamp 1626908933
transform 1 0 30336 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_693
timestamp 1626908933
transform 1 0 30336 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_124
timestamp 1626908933
transform 1 0 29952 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_693
timestamp 1626908933
transform 1 0 29952 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_570
timestamp 1626908933
transform 1 0 31104 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_202
timestamp 1626908933
transform 1 0 31104 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_676
timestamp 1626908933
transform 1 0 31296 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_107
timestamp 1626908933
transform 1 0 31296 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_579
timestamp 1626908933
transform 1 0 31104 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_211
timestamp 1626908933
transform 1 0 31104 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_677
timestamp 1626908933
transform 1 0 31296 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_108
timestamp 1626908933
transform 1 0 31296 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_668
timestamp 1626908933
transform 1 0 31680 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_98
timestamp 1626908933
transform 1 0 31680 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_669
timestamp 1626908933
transform 1 0 31680 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_99
timestamp 1626908933
transform 1 0 31680 0 1 2664
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_301
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_13
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_282
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_12
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_282
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_12
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_282
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_12
timestamp 1626908933
transform 1 0 32600 0 1 3330
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_466
timestamp 1626908933
transform 1 0 32448 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_207
timestamp 1626908933
transform 1 0 32448 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_981
timestamp 1626908933
transform 1 0 32448 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_351
timestamp 1626908933
transform 1 0 32448 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_76
timestamp 1626908933
transform 1 0 32544 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_645
timestamp 1626908933
transform 1 0 32544 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_75
timestamp 1626908933
transform 1 0 32544 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_644
timestamp 1626908933
transform 1 0 32544 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_639
timestamp 1626908933
transform 1 0 32928 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_69
timestamp 1626908933
transform 1 0 32928 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_640
timestamp 1626908933
transform 1 0 32928 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_70
timestamp 1626908933
transform 1 0 32928 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_350
timestamp 1626908933
transform 1 0 33696 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_980
timestamp 1626908933
transform 1 0 33696 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_330
timestamp 1626908933
transform 1 0 33696 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_960
timestamp 1626908933
transform 1 0 33696 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_40
timestamp 1626908933
transform 1 0 34176 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_610
timestamp 1626908933
transform 1 0 34176 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_43
timestamp 1626908933
transform 1 0 33792 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_612
timestamp 1626908933
transform 1 0 33792 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_39
timestamp 1626908933
transform 1 0 34176 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_609
timestamp 1626908933
transform 1 0 34176 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_42
timestamp 1626908933
transform 1 0 33792 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_611
timestamp 1626908933
transform 1 0 33792 0 -1 3996
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_418
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_148
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_418
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_148
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_418
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_148
timestamp 1626908933
transform 1 0 34600 0 1 2664
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_582
timestamp 1626908933
transform 1 0 34944 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_12
timestamp 1626908933
transform 1 0 34944 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_631
timestamp 1626908933
transform 1 0 35424 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_263
timestamp 1626908933
transform 1 0 35424 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_582
timestamp 1626908933
transform 1 0 35040 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_13
timestamp 1626908933
transform 1 0 35040 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_473
timestamp 1626908933
transform 1 0 34944 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_214
timestamp 1626908933
transform 1 0 34944 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1092
timestamp 1626908933
transform 1 0 35616 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_462
timestamp 1626908933
transform 1 0 35616 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_465
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_206
timestamp 1626908933
transform 1 0 288 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1137
timestamp 1626908933
transform 1 0 480 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_568
timestamp 1626908933
transform 1 0 480 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_3
timestamp 1626908933
transform 1 0 864 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_23
timestamp 1626908933
transform 1 0 864 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_959
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_329
timestamp 1626908933
transform 1 0 384 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_958
timestamp 1626908933
transform 1 0 1344 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_328
timestamp 1626908933
transform 1 0 1344 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1363
timestamp 1626908933
transform 1 0 1296 0 1 3589
box -29 -23 29 23
use L1M1_PR  L1M1_PR_575
timestamp 1626908933
transform 1 0 1296 0 1 3589
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1271
timestamp 1626908933
transform 1 0 1296 0 1 3589
box -32 -32 32 32
use M1M2_PR  M1M2_PR_503
timestamp 1626908933
transform 1 0 1296 0 1 3589
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1135
timestamp 1626908933
transform 1 0 1440 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_565
timestamp 1626908933
transform 1 0 1440 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_957
timestamp 1626908933
transform 1 0 2208 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_327
timestamp 1626908933
transform 1 0 2208 0 1 3996
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1369
timestamp 1626908933
transform 1 0 1584 0 1 3737
box -29 -23 29 23
use L1M1_PR  L1M1_PR_581
timestamp 1626908933
transform 1 0 1584 0 1 3737
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1277
timestamp 1626908933
transform 1 0 2064 0 1 3737
box -32 -32 32 32
use M1M2_PR  M1M2_PR_509
timestamp 1626908933
transform 1 0 2064 0 1 3737
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_267
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_537
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_267
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_537
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_267
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_537
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_284
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_572
timestamp 1626908933
transform 1 0 2600 0 1 3996
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_549
timestamp 1626908933
transform 1 0 2688 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1119
timestamp 1626908933
transform 1 0 2688 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_547
timestamp 1626908933
transform 1 0 2304 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1116
timestamp 1626908933
transform 1 0 2304 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_956
timestamp 1626908933
transform 1 0 3456 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_326
timestamp 1626908933
transform 1 0 3456 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1099
timestamp 1626908933
transform 1 0 3552 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_530
timestamp 1626908933
transform 1 0 3552 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_955
timestamp 1626908933
transform 1 0 3936 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_325
timestamp 1626908933
transform 1 0 3936 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1110
timestamp 1626908933
transform 1 0 4032 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_540
timestamp 1626908933
transform 1 0 4032 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_632
timestamp 1626908933
transform 1 0 4800 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_264
timestamp 1626908933
transform 1 0 4800 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_464
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_205
timestamp 1626908933
transform 1 0 4992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_569
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_201
timestamp 1626908933
transform 1 0 5088 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1096
timestamp 1626908933
transform 1 0 5280 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_526
timestamp 1626908933
transform 1 0 5280 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_324
timestamp 1626908933
transform 1 0 6048 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_954
timestamp 1626908933
transform 1 0 6048 0 1 3996
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_556
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_268
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_522
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_252
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_522
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_252
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_522
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_252
timestamp 1626908933
transform 1 0 6600 0 1 3996
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_953
timestamp 1626908933
transform 1 0 6528 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_323
timestamp 1626908933
transform 1 0 6528 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_512
timestamp 1626908933
transform 1 0 6624 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1082
timestamp 1626908933
transform 1 0 6624 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_501
timestamp 1626908933
transform 1 0 6144 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1070
timestamp 1626908933
transform 1 0 6144 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_952
timestamp 1626908933
transform 1 0 7392 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_322
timestamp 1626908933
transform 1 0 7392 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1057
timestamp 1626908933
transform 1 0 7488 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_488
timestamp 1626908933
transform 1 0 7488 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1064
timestamp 1626908933
transform 1 0 7872 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_494
timestamp 1626908933
transform 1 0 7872 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_951
timestamp 1626908933
transform 1 0 8640 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_321
timestamp 1626908933
transform 1 0 8640 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1043
timestamp 1626908933
transform 1 0 8736 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_474
timestamp 1626908933
transform 1 0 8736 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1050
timestamp 1626908933
transform 1 0 9120 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_480
timestamp 1626908933
transform 1 0 9120 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_204
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_463
timestamp 1626908933
transform 1 0 9984 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_465
timestamp 1626908933
transform 1 0 9888 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1095
timestamp 1626908933
transform 1 0 9888 0 1 3996
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_540
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_252
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_237
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_507
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_237
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_507
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_237
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_507
timestamp 1626908933
transform 1 0 10600 0 1 3996
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_467
timestamp 1626908933
transform 1 0 10464 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1037
timestamp 1626908933
transform 1 0 10464 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_450
timestamp 1626908933
transform 1 0 10080 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1019
timestamp 1626908933
transform 1 0 10080 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_950
timestamp 1626908933
transform 1 0 11232 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_320
timestamp 1626908933
transform 1 0 11232 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_998
timestamp 1626908933
transform 1 0 11328 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_429
timestamp 1626908933
transform 1 0 11328 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1016
timestamp 1626908933
transform 1 0 11712 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_446
timestamp 1626908933
transform 1 0 11712 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_978
timestamp 1626908933
transform 1 0 12480 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_409
timestamp 1626908933
transform 1 0 12480 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_949
timestamp 1626908933
transform 1 0 12864 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_319
timestamp 1626908933
transform 1 0 12864 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1003
timestamp 1626908933
transform 1 0 12960 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_433
timestamp 1626908933
transform 1 0 12960 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_948
timestamp 1626908933
transform 1 0 13728 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_318
timestamp 1626908933
transform 1 0 13728 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_950
timestamp 1626908933
transform 1 0 13824 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_381
timestamp 1626908933
transform 1 0 13824 0 1 3996
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_524
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_236
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_222
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_492
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_222
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_492
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_222
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_492
timestamp 1626908933
transform 1 0 14600 0 1 3996
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_203
timestamp 1626908933
transform 1 0 14976 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_462
timestamp 1626908933
transform 1 0 14976 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_419
timestamp 1626908933
transform 1 0 14208 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_989
timestamp 1626908933
transform 1 0 14208 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_947
timestamp 1626908933
transform 1 0 15072 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_317
timestamp 1626908933
transform 1 0 15072 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_931
timestamp 1626908933
transform 1 0 15168 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_362
timestamp 1626908933
transform 1 0 15168 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_969
timestamp 1626908933
transform 1 0 15552 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_399
timestamp 1626908933
transform 1 0 15552 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_943
timestamp 1626908933
transform 1 0 16896 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_373
timestamp 1626908933
transform 1 0 16896 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_568
timestamp 1626908933
transform 1 0 16320 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_200
timestamp 1626908933
transform 1 0 16320 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_906
timestamp 1626908933
transform 1 0 16512 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_337
timestamp 1626908933
transform 1 0 16512 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_946
timestamp 1626908933
transform 1 0 17664 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_316
timestamp 1626908933
transform 1 0 17664 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_881
timestamp 1626908933
transform 1 0 17760 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_312
timestamp 1626908933
transform 1 0 17760 0 1 3996
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_508
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_220
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_207
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_477
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_207
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_477
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_207
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_477
timestamp 1626908933
transform 1 0 18600 0 1 3996
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_350
timestamp 1626908933
transform 1 0 18144 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_920
timestamp 1626908933
transform 1 0 18144 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_945
timestamp 1626908933
transform 1 0 19104 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_315
timestamp 1626908933
transform 1 0 19104 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_567
timestamp 1626908933
transform 1 0 18912 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_199
timestamp 1626908933
transform 1 0 18912 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_898
timestamp 1626908933
transform 1 0 19200 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_328
timestamp 1626908933
transform 1 0 19200 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_876
timestamp 1626908933
transform 1 0 20064 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_306
timestamp 1626908933
transform 1 0 20064 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_461
timestamp 1626908933
transform 1 0 19968 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_202
timestamp 1626908933
transform 1 0 19968 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_566
timestamp 1626908933
transform 1 0 20832 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_198
timestamp 1626908933
transform 1 0 20832 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_827
timestamp 1626908933
transform 1 0 21024 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_258
timestamp 1626908933
transform 1 0 21024 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_850
timestamp 1626908933
transform 1 0 21408 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_280
timestamp 1626908933
transform 1 0 21408 0 1 3996
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_492
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_204
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_462
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_192
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_462
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_192
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_462
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_192
timestamp 1626908933
transform 1 0 22600 0 1 3996
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_944
timestamp 1626908933
transform 1 0 22176 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_314
timestamp 1626908933
transform 1 0 22176 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_239
timestamp 1626908933
transform 1 0 22272 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_808
timestamp 1626908933
transform 1 0 22272 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_828
timestamp 1626908933
transform 1 0 22656 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_258
timestamp 1626908933
transform 1 0 22656 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_793
timestamp 1626908933
transform 1 0 23424 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_224
timestamp 1626908933
transform 1 0 23424 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_943
timestamp 1626908933
transform 1 0 23808 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_313
timestamp 1626908933
transform 1 0 23808 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_805
timestamp 1626908933
transform 1 0 23904 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_235
timestamp 1626908933
transform 1 0 23904 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_565
timestamp 1626908933
transform 1 0 25056 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_197
timestamp 1626908933
transform 1 0 25056 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_460
timestamp 1626908933
transform 1 0 24960 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_201
timestamp 1626908933
transform 1 0 24960 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_633
timestamp 1626908933
transform 1 0 24672 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_265
timestamp 1626908933
transform 1 0 24672 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1096
timestamp 1626908933
transform 1 0 24864 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_466
timestamp 1626908933
transform 1 0 24864 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_784
timestamp 1626908933
transform 1 0 25248 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_214
timestamp 1626908933
transform 1 0 25248 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_756
timestamp 1626908933
transform 1 0 26016 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_187
timestamp 1626908933
transform 1 0 26016 0 1 3996
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_476
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_188
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_447
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_177
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_447
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_177
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_447
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_177
timestamp 1626908933
transform 1 0 26600 0 1 3996
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_942
timestamp 1626908933
transform 1 0 26400 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_312
timestamp 1626908933
transform 1 0 26400 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_192
timestamp 1626908933
transform 1 0 26496 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_762
timestamp 1626908933
transform 1 0 26496 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_740
timestamp 1626908933
transform 1 0 27840 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_170
timestamp 1626908933
transform 1 0 27840 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_564
timestamp 1626908933
transform 1 0 27264 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_196
timestamp 1626908933
transform 1 0 27264 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_735
timestamp 1626908933
transform 1 0 27456 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_166
timestamp 1626908933
transform 1 0 27456 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_719
timestamp 1626908933
transform 1 0 28608 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_150
timestamp 1626908933
transform 1 0 28608 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_941
timestamp 1626908933
transform 1 0 28992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_311
timestamp 1626908933
transform 1 0 28992 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_716
timestamp 1626908933
transform 1 0 29088 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_146
timestamp 1626908933
transform 1 0 29088 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1097
timestamp 1626908933
transform 1 0 29856 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_467
timestamp 1626908933
transform 1 0 29856 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_310
timestamp 1626908933
transform 1 0 30240 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_940
timestamp 1626908933
transform 1 0 30240 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_200
timestamp 1626908933
transform 1 0 29952 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_459
timestamp 1626908933
transform 1 0 29952 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_195
timestamp 1626908933
transform 1 0 30048 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_563
timestamp 1626908933
transform 1 0 30048 0 1 3996
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_162
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_432
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_162
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_432
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_162
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_432
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_172
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_460
timestamp 1626908933
transform 1 0 30600 0 1 3996
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_122
timestamp 1626908933
transform 1 0 30336 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_692
timestamp 1626908933
transform 1 0 30336 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_562
timestamp 1626908933
transform 1 0 31104 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_194
timestamp 1626908933
transform 1 0 31104 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_675
timestamp 1626908933
transform 1 0 31296 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_106
timestamp 1626908933
transform 1 0 31296 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_667
timestamp 1626908933
transform 1 0 31680 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_97
timestamp 1626908933
transform 1 0 31680 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_939
timestamp 1626908933
transform 1 0 32448 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_309
timestamp 1626908933
transform 1 0 32448 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_643
timestamp 1626908933
transform 1 0 32544 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_74
timestamp 1626908933
transform 1 0 32544 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_638
timestamp 1626908933
transform 1 0 32928 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_68
timestamp 1626908933
transform 1 0 32928 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_938
timestamp 1626908933
transform 1 0 33696 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_308
timestamp 1626908933
transform 1 0 33696 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_610
timestamp 1626908933
transform 1 0 33792 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_41
timestamp 1626908933
transform 1 0 33792 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_608
timestamp 1626908933
transform 1 0 34176 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_38
timestamp 1626908933
transform 1 0 34176 0 1 3996
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_417
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_147
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_417
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_147
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_417
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_147
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_156
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_444
timestamp 1626908933
transform 1 0 34600 0 1 3996
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_199
timestamp 1626908933
transform 1 0 34944 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_458
timestamp 1626908933
transform 1 0 34944 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_12
timestamp 1626908933
transform 1 0 35040 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_581
timestamp 1626908933
transform 1 0 35040 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_266
timestamp 1626908933
transform 1 0 35424 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_634
timestamp 1626908933
transform 1 0 35424 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_468
timestamp 1626908933
transform 1 0 35616 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1098
timestamp 1626908933
transform 1 0 35616 0 1 3996
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1525
timestamp 1626908933
transform 1 0 48 0 1 4847
box -32 -32 32 32
use M1M2_PR  M1M2_PR_757
timestamp 1626908933
transform 1 0 48 0 1 4847
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1099
timestamp 1626908933
transform 1 0 288 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_469
timestamp 1626908933
transform 1 0 288 0 -1 5328
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_428
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_140
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_131
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_401
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_131
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_401
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_131
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_401
timestamp 1626908933
transform 1 0 600 0 1 4662
box -200 -49 200 49
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_21
timestamp 1626908933
transform 1 0 384 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_1
timestamp 1626908933
transform 1 0 384 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_561
timestamp 1626908933
transform 1 0 864 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1130
timestamp 1626908933
transform 1 0 864 0 -1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_342
timestamp 1626908933
transform 1 0 1008 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_763
timestamp 1626908933
transform 1 0 912 0 1 4329
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1110
timestamp 1626908933
transform 1 0 1008 0 1 4551
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1531
timestamp 1626908933
transform 1 0 912 0 1 4329
box -32 -32 32 32
use L1M1_PR  L1M1_PR_414
timestamp 1626908933
transform 1 0 1008 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_785
timestamp 1626908933
transform 1 0 912 0 1 4329
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1202
timestamp 1626908933
transform 1 0 1008 0 1 4551
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1573
timestamp 1626908933
transform 1 0 912 0 1 4329
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_193
timestamp 1626908933
transform 1 0 1248 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_561
timestamp 1626908933
transform 1 0 1248 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1134
timestamp 1626908933
transform 1 0 1440 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_564
timestamp 1626908933
transform 1 0 1440 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_560
timestamp 1626908933
transform 1 0 2208 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_192
timestamp 1626908933
transform 1 0 2208 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1100
timestamp 1626908933
transform 1 0 2400 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_470
timestamp 1626908933
transform 1 0 2400 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_457
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_198
timestamp 1626908933
transform 1 0 2496 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_937
timestamp 1626908933
transform 1 0 2592 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_307
timestamp 1626908933
transform 1 0 2592 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1118
timestamp 1626908933
transform 1 0 2688 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_548
timestamp 1626908933
transform 1 0 2688 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_936
timestamp 1626908933
transform 1 0 3456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_306
timestamp 1626908933
transform 1 0 3456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1098
timestamp 1626908933
transform 1 0 3552 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_529
timestamp 1626908933
transform 1 0 3552 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_935
timestamp 1626908933
transform 1 0 3936 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_305
timestamp 1626908933
transform 1 0 3936 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1109
timestamp 1626908933
transform 1 0 4032 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_539
timestamp 1626908933
transform 1 0 4032 0 -1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1329
timestamp 1626908933
transform 1 0 4080 0 1 4403
box -32 -32 32 32
use M1M2_PR  M1M2_PR_561
timestamp 1626908933
transform 1 0 4080 0 1 4403
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_124
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_412
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_116
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_386
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_116
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_386
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_116
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_386
timestamp 1626908933
transform 1 0 4600 0 1 4662
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_304
timestamp 1626908933
transform 1 0 4800 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_934
timestamp 1626908933
transform 1 0 4800 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_519
timestamp 1626908933
transform 1 0 4896 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1088
timestamp 1626908933
transform 1 0 4896 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1095
timestamp 1626908933
transform 1 0 5280 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_525
timestamp 1626908933
transform 1 0 5280 0 -1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1516
timestamp 1626908933
transform 1 0 5424 0 1 4847
box -32 -32 32 32
use M1M2_PR  M1M2_PR_748
timestamp 1626908933
transform 1 0 5424 0 1 4847
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_933
timestamp 1626908933
transform 1 0 6048 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_303
timestamp 1626908933
transform 1 0 6048 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1069
timestamp 1626908933
transform 1 0 6144 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_500
timestamp 1626908933
transform 1 0 6144 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1081
timestamp 1626908933
transform 1 0 6624 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_511
timestamp 1626908933
transform 1 0 6624 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_932
timestamp 1626908933
transform 1 0 6528 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_302
timestamp 1626908933
transform 1 0 6528 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_931
timestamp 1626908933
transform 1 0 7776 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_301
timestamp 1626908933
transform 1 0 7776 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1101
timestamp 1626908933
transform 1 0 7392 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_471
timestamp 1626908933
transform 1 0 7392 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_559
timestamp 1626908933
transform 1 0 7584 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_191
timestamp 1626908933
transform 1 0 7584 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_456
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_197
timestamp 1626908933
transform 1 0 7488 0 -1 5328
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_108
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_396
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_101
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_371
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_101
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_371
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_101
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_371
timestamp 1626908933
transform 1 0 8600 0 1 4662
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_493
timestamp 1626908933
transform 1 0 7872 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1063
timestamp 1626908933
transform 1 0 7872 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1042
timestamp 1626908933
transform 1 0 8736 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_473
timestamp 1626908933
transform 1 0 8736 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1049
timestamp 1626908933
transform 1 0 9120 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_479
timestamp 1626908933
transform 1 0 9120 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_930
timestamp 1626908933
transform 1 0 8640 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_300
timestamp 1626908933
transform 1 0 8640 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1025
timestamp 1626908933
transform 1 0 9888 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_456
timestamp 1626908933
transform 1 0 9888 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1036
timestamp 1626908933
transform 1 0 10464 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_466
timestamp 1626908933
transform 1 0 10464 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_558
timestamp 1626908933
transform 1 0 10272 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_190
timestamp 1626908933
transform 1 0 10272 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_997
timestamp 1626908933
transform 1 0 11328 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_428
timestamp 1626908933
transform 1 0 11328 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_929
timestamp 1626908933
transform 1 0 11232 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_299
timestamp 1626908933
transform 1 0 11232 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1015
timestamp 1626908933
transform 1 0 11712 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_445
timestamp 1626908933
transform 1 0 11712 0 -1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1327
timestamp 1626908933
transform 1 0 11760 0 1 4255
box -32 -32 32 32
use M1M2_PR  M1M2_PR_559
timestamp 1626908933
transform 1 0 11760 0 1 4255
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_356
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_86
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_356
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_86
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_356
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_86
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_380
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_92
timestamp 1626908933
transform 1 0 12600 0 1 4662
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_969
timestamp 1626908933
transform 1 0 12576 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_400
timestamp 1626908933
transform 1 0 12576 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_455
timestamp 1626908933
transform 1 0 12480 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_196
timestamp 1626908933
transform 1 0 12480 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1002
timestamp 1626908933
transform 1 0 12960 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_432
timestamp 1626908933
transform 1 0 12960 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_949
timestamp 1626908933
transform 1 0 13920 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_380
timestamp 1626908933
transform 1 0 13920 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_557
timestamp 1626908933
transform 1 0 13728 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_189
timestamp 1626908933
transform 1 0 13728 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_988
timestamp 1626908933
transform 1 0 14304 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_418
timestamp 1626908933
transform 1 0 14304 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_930
timestamp 1626908933
transform 1 0 15168 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_361
timestamp 1626908933
transform 1 0 15168 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_928
timestamp 1626908933
transform 1 0 15072 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_298
timestamp 1626908933
transform 1 0 15072 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_968
timestamp 1626908933
transform 1 0 15552 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_398
timestamp 1626908933
transform 1 0 15552 0 -1 5328
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_76
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_364
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_71
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_341
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_71
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_341
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_71
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_341
timestamp 1626908933
transform 1 0 16600 0 1 4662
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_336
timestamp 1626908933
transform 1 0 16320 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_905
timestamp 1626908933
transform 1 0 16320 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_372
timestamp 1626908933
transform 1 0 16704 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_942
timestamp 1626908933
transform 1 0 16704 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_454
timestamp 1626908933
transform 1 0 17472 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_195
timestamp 1626908933
transform 1 0 17472 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_880
timestamp 1626908933
transform 1 0 17760 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_311
timestamp 1626908933
transform 1 0 17760 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_556
timestamp 1626908933
transform 1 0 17568 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_188
timestamp 1626908933
transform 1 0 17568 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_919
timestamp 1626908933
transform 1 0 18144 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_349
timestamp 1626908933
transform 1 0 18144 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_858
timestamp 1626908933
transform 1 0 18912 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_289
timestamp 1626908933
transform 1 0 18912 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_927
timestamp 1626908933
transform 1 0 19296 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_297
timestamp 1626908933
transform 1 0 19296 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_897
timestamp 1626908933
transform 1 0 19392 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_327
timestamp 1626908933
transform 1 0 19392 0 -1 5328
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_326
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_56
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_326
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_56
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_326
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_56
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_348
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_60
timestamp 1626908933
transform 1 0 20600 0 1 4662
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_555
timestamp 1626908933
transform 1 0 20160 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_187
timestamp 1626908933
transform 1 0 20160 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_273
timestamp 1626908933
transform 1 0 20352 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_842
timestamp 1626908933
transform 1 0 20352 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_864
timestamp 1626908933
transform 1 0 20736 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_294
timestamp 1626908933
transform 1 0 20736 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_554
timestamp 1626908933
transform 1 0 21504 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_186
timestamp 1626908933
transform 1 0 21504 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_840
timestamp 1626908933
transform 1 0 21696 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_270
timestamp 1626908933
transform 1 0 21696 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_827
timestamp 1626908933
transform 1 0 22656 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_257
timestamp 1626908933
transform 1 0 22656 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_926
timestamp 1626908933
transform 1 0 22560 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_296
timestamp 1626908933
transform 1 0 22560 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_453
timestamp 1626908933
transform 1 0 22464 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_194
timestamp 1626908933
transform 1 0 22464 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_792
timestamp 1626908933
transform 1 0 23424 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_223
timestamp 1626908933
transform 1 0 23424 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_925
timestamp 1626908933
transform 1 0 23808 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_295
timestamp 1626908933
transform 1 0 23808 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_804
timestamp 1626908933
transform 1 0 23904 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_234
timestamp 1626908933
transform 1 0 23904 0 -1 5328
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_311
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_41
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_311
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_41
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_311
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_41
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_332
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_44
timestamp 1626908933
transform 1 0 24600 0 1 4662
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_553
timestamp 1626908933
transform 1 0 24672 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_185
timestamp 1626908933
transform 1 0 24672 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_203
timestamp 1626908933
transform 1 0 24864 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_772
timestamp 1626908933
transform 1 0 24864 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_783
timestamp 1626908933
transform 1 0 25248 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_213
timestamp 1626908933
transform 1 0 25248 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_755
timestamp 1626908933
transform 1 0 26016 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_186
timestamp 1626908933
transform 1 0 26016 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_761
timestamp 1626908933
transform 1 0 26496 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_191
timestamp 1626908933
transform 1 0 26496 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_924
timestamp 1626908933
transform 1 0 26400 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_294
timestamp 1626908933
transform 1 0 26400 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_184
timestamp 1626908933
transform 1 0 27552 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_552
timestamp 1626908933
transform 1 0 27552 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_193
timestamp 1626908933
transform 1 0 27456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_452
timestamp 1626908933
transform 1 0 27456 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_293
timestamp 1626908933
transform 1 0 27264 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_472
timestamp 1626908933
transform 1 0 27360 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_923
timestamp 1626908933
transform 1 0 27264 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1102
timestamp 1626908933
transform 1 0 27360 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_292
timestamp 1626908933
transform 1 0 27744 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_922
timestamp 1626908933
transform 1 0 27744 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_169
timestamp 1626908933
transform 1 0 27840 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_739
timestamp 1626908933
transform 1 0 27840 0 -1 5328
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_28
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_316
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_26
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_296
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_26
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_296
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_26
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_296
timestamp 1626908933
transform 1 0 28600 0 1 4662
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_149
timestamp 1626908933
transform 1 0 28608 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_718
timestamp 1626908933
transform 1 0 28608 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_921
timestamp 1626908933
transform 1 0 28992 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_291
timestamp 1626908933
transform 1 0 28992 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_715
timestamp 1626908933
transform 1 0 29088 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_145
timestamp 1626908933
transform 1 0 29088 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_920
timestamp 1626908933
transform 1 0 29856 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_290
timestamp 1626908933
transform 1 0 29856 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_692
timestamp 1626908933
transform 1 0 29952 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_123
timestamp 1626908933
transform 1 0 29952 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_691
timestamp 1626908933
transform 1 0 30336 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_121
timestamp 1626908933
transform 1 0 30336 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_551
timestamp 1626908933
transform 1 0 31104 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_183
timestamp 1626908933
transform 1 0 31104 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_674
timestamp 1626908933
transform 1 0 31296 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_105
timestamp 1626908933
transform 1 0 31296 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_666
timestamp 1626908933
transform 1 0 31680 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_96
timestamp 1626908933
transform 1 0 31680 0 -1 5328
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_281
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_11
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_281
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_11
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_281
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_11
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_300
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_12
timestamp 1626908933
transform 1 0 32600 0 1 4662
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_451
timestamp 1626908933
transform 1 0 32448 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_192
timestamp 1626908933
transform 1 0 32448 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_73
timestamp 1626908933
transform 1 0 32544 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_642
timestamp 1626908933
transform 1 0 32544 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_637
timestamp 1626908933
transform 1 0 32928 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_67
timestamp 1626908933
transform 1 0 32928 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_919
timestamp 1626908933
transform 1 0 33696 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_289
timestamp 1626908933
transform 1 0 33696 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_609
timestamp 1626908933
transform 1 0 33792 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_40
timestamp 1626908933
transform 1 0 33792 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_607
timestamp 1626908933
transform 1 0 34176 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_37
timestamp 1626908933
transform 1 0 34176 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_11
timestamp 1626908933
transform 1 0 34944 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_581
timestamp 1626908933
transform 1 0 34944 0 -1 5328
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1503
timestamp 1626908933
transform 1 0 48 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_735
timestamp 1626908933
transform 1 0 48 0 1 5513
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1193
timestamp 1626908933
transform 1 0 144 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_405
timestamp 1626908933
transform 1 0 144 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_450
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_191
timestamp 1626908933
transform 1 0 288 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1129
timestamp 1626908933
transform 1 0 864 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_560
timestamp 1626908933
transform 1 0 864 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_2
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_22
timestamp 1626908933
transform 1 0 384 0 1 5328
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1191
timestamp 1626908933
transform 1 0 528 0 1 5217
box -29 -23 29 23
use L1M1_PR  L1M1_PR_403
timestamp 1626908933
transform 1 0 528 0 1 5217
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_550
timestamp 1626908933
transform 1 0 1248 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_182
timestamp 1626908933
transform 1 0 1248 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1133
timestamp 1626908933
transform 1 0 1440 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_563
timestamp 1626908933
transform 1 0 1440 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1117
timestamp 1626908933
transform 1 0 2208 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_547
timestamp 1626908933
transform 1 0 2208 0 1 5328
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_283
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_571
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_266
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_536
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_266
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_536
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_266
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_536
timestamp 1626908933
transform 1 0 2600 0 1 5328
box -200 -49 200 49
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_101
timestamp 1626908933
transform 1 0 2976 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_46
timestamp 1626908933
transform 1 0 2976 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_45
timestamp 1626908933
transform 1 0 3456 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_100
timestamp 1626908933
transform 1 0 3456 0 1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_918
timestamp 1626908933
transform 1 0 3936 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_288
timestamp 1626908933
transform 1 0 3936 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1108
timestamp 1626908933
transform 1 0 4032 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_538
timestamp 1626908933
transform 1 0 4032 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_449
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_190
timestamp 1626908933
transform 1 0 4992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1103
timestamp 1626908933
transform 1 0 4896 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_917
timestamp 1626908933
transform 1 0 4800 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_473
timestamp 1626908933
transform 1 0 4896 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_287
timestamp 1626908933
transform 1 0 4800 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1094
timestamp 1626908933
transform 1 0 5280 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_524
timestamp 1626908933
transform 1 0 5280 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_549
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_181
timestamp 1626908933
transform 1 0 5088 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_286
timestamp 1626908933
transform 1 0 6048 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_916
timestamp 1626908933
transform 1 0 6048 0 1 5328
box -38 -49 134 715
use M1M2_PR  M1M2_PR_734
timestamp 1626908933
transform 1 0 6000 0 1 5513
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1502
timestamp 1626908933
transform 1 0 6000 0 1 5513
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_555
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_267
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_521
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_251
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_521
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_251
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_521
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_251
timestamp 1626908933
transform 1 0 6600 0 1 5328
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_915
timestamp 1626908933
transform 1 0 6528 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_285
timestamp 1626908933
transform 1 0 6528 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_510
timestamp 1626908933
transform 1 0 6624 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1080
timestamp 1626908933
transform 1 0 6624 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_499
timestamp 1626908933
transform 1 0 6144 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1068
timestamp 1626908933
transform 1 0 6144 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1056
timestamp 1626908933
transform 1 0 7488 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_487
timestamp 1626908933
transform 1 0 7488 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_914
timestamp 1626908933
transform 1 0 7392 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_284
timestamp 1626908933
transform 1 0 7392 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1062
timestamp 1626908933
transform 1 0 7872 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_492
timestamp 1626908933
transform 1 0 7872 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1041
timestamp 1626908933
transform 1 0 8736 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_472
timestamp 1626908933
transform 1 0 8736 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1048
timestamp 1626908933
transform 1 0 9120 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_478
timestamp 1626908933
transform 1 0 9120 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_913
timestamp 1626908933
transform 1 0 8640 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_283
timestamp 1626908933
transform 1 0 8640 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_189
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_448
timestamp 1626908933
transform 1 0 9984 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_474
timestamp 1626908933
transform 1 0 9888 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1104
timestamp 1626908933
transform 1 0 9888 0 1 5328
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_236
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_506
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_236
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_506
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_236
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_506
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_251
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_539
timestamp 1626908933
transform 1 0 10600 0 1 5328
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_465
timestamp 1626908933
transform 1 0 10464 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1035
timestamp 1626908933
transform 1 0 10464 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_449
timestamp 1626908933
transform 1 0 10080 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1018
timestamp 1626908933
transform 1 0 10080 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_996
timestamp 1626908933
transform 1 0 11328 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_427
timestamp 1626908933
transform 1 0 11328 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_912
timestamp 1626908933
transform 1 0 11232 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_282
timestamp 1626908933
transform 1 0 11232 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1014
timestamp 1626908933
transform 1 0 11712 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_444
timestamp 1626908933
transform 1 0 11712 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_977
timestamp 1626908933
transform 1 0 12480 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_408
timestamp 1626908933
transform 1 0 12480 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_911
timestamp 1626908933
transform 1 0 12864 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_281
timestamp 1626908933
transform 1 0 12864 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1001
timestamp 1626908933
transform 1 0 12960 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_431
timestamp 1626908933
transform 1 0 12960 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_910
timestamp 1626908933
transform 1 0 13728 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_280
timestamp 1626908933
transform 1 0 13728 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_948
timestamp 1626908933
transform 1 0 13824 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_379
timestamp 1626908933
transform 1 0 13824 0 1 5328
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_523
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_235
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_221
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_491
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_221
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_491
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_221
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_491
timestamp 1626908933
transform 1 0 14600 0 1 5328
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_188
timestamp 1626908933
transform 1 0 14976 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_447
timestamp 1626908933
transform 1 0 14976 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_417
timestamp 1626908933
transform 1 0 14208 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_987
timestamp 1626908933
transform 1 0 14208 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_929
timestamp 1626908933
transform 1 0 15168 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_360
timestamp 1626908933
transform 1 0 15168 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_909
timestamp 1626908933
transform 1 0 15072 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_279
timestamp 1626908933
transform 1 0 15072 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_967
timestamp 1626908933
transform 1 0 15552 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_397
timestamp 1626908933
transform 1 0 15552 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_941
timestamp 1626908933
transform 1 0 16896 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_371
timestamp 1626908933
transform 1 0 16896 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_548
timestamp 1626908933
transform 1 0 16320 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_180
timestamp 1626908933
transform 1 0 16320 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_904
timestamp 1626908933
transform 1 0 16512 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_335
timestamp 1626908933
transform 1 0 16512 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_879
timestamp 1626908933
transform 1 0 17760 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_310
timestamp 1626908933
transform 1 0 17760 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_908
timestamp 1626908933
transform 1 0 17664 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_278
timestamp 1626908933
transform 1 0 17664 0 1 5328
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_507
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_219
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_206
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_476
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_206
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_476
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_206
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_476
timestamp 1626908933
transform 1 0 18600 0 1 5328
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_348
timestamp 1626908933
transform 1 0 18144 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_918
timestamp 1626908933
transform 1 0 18144 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_907
timestamp 1626908933
transform 1 0 19104 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_277
timestamp 1626908933
transform 1 0 19104 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_547
timestamp 1626908933
transform 1 0 18912 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_179
timestamp 1626908933
transform 1 0 18912 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_896
timestamp 1626908933
transform 1 0 19200 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_326
timestamp 1626908933
transform 1 0 19200 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_875
timestamp 1626908933
transform 1 0 20064 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_305
timestamp 1626908933
transform 1 0 20064 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_446
timestamp 1626908933
transform 1 0 19968 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_187
timestamp 1626908933
transform 1 0 19968 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_826
timestamp 1626908933
transform 1 0 21024 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_257
timestamp 1626908933
transform 1 0 21024 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_546
timestamp 1626908933
transform 1 0 20832 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_178
timestamp 1626908933
transform 1 0 20832 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_849
timestamp 1626908933
transform 1 0 21408 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_279
timestamp 1626908933
transform 1 0 21408 0 1 5328
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_491
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_203
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_461
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_191
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_461
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_191
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_461
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_191
timestamp 1626908933
transform 1 0 22600 0 1 5328
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_906
timestamp 1626908933
transform 1 0 22176 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_276
timestamp 1626908933
transform 1 0 22176 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_238
timestamp 1626908933
transform 1 0 22272 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_807
timestamp 1626908933
transform 1 0 22272 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_826
timestamp 1626908933
transform 1 0 22656 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_256
timestamp 1626908933
transform 1 0 22656 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_791
timestamp 1626908933
transform 1 0 23424 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_222
timestamp 1626908933
transform 1 0 23424 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_905
timestamp 1626908933
transform 1 0 23808 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_275
timestamp 1626908933
transform 1 0 23808 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_803
timestamp 1626908933
transform 1 0 23904 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_233
timestamp 1626908933
transform 1 0 23904 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_545
timestamp 1626908933
transform 1 0 25056 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_177
timestamp 1626908933
transform 1 0 25056 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_445
timestamp 1626908933
transform 1 0 24960 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_186
timestamp 1626908933
transform 1 0 24960 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_635
timestamp 1626908933
transform 1 0 24672 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_267
timestamp 1626908933
transform 1 0 24672 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1105
timestamp 1626908933
transform 1 0 24864 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_475
timestamp 1626908933
transform 1 0 24864 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_782
timestamp 1626908933
transform 1 0 25248 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_212
timestamp 1626908933
transform 1 0 25248 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_754
timestamp 1626908933
transform 1 0 26016 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_185
timestamp 1626908933
transform 1 0 26016 0 1 5328
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_475
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_187
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_446
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_176
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_446
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_176
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_446
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_176
timestamp 1626908933
transform 1 0 26600 0 1 5328
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_904
timestamp 1626908933
transform 1 0 26400 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_274
timestamp 1626908933
transform 1 0 26400 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_190
timestamp 1626908933
transform 1 0 26496 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_760
timestamp 1626908933
transform 1 0 26496 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_738
timestamp 1626908933
transform 1 0 27840 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_168
timestamp 1626908933
transform 1 0 27840 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_734
timestamp 1626908933
transform 1 0 27456 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_165
timestamp 1626908933
transform 1 0 27456 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_544
timestamp 1626908933
transform 1 0 27264 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_176
timestamp 1626908933
transform 1 0 27264 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_717
timestamp 1626908933
transform 1 0 28608 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_148
timestamp 1626908933
transform 1 0 28608 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_903
timestamp 1626908933
transform 1 0 28992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_273
timestamp 1626908933
transform 1 0 28992 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_714
timestamp 1626908933
transform 1 0 29088 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_144
timestamp 1626908933
transform 1 0 29088 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1106
timestamp 1626908933
transform 1 0 29856 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_476
timestamp 1626908933
transform 1 0 29856 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_272
timestamp 1626908933
transform 1 0 30240 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_902
timestamp 1626908933
transform 1 0 30240 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_185
timestamp 1626908933
transform 1 0 29952 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_444
timestamp 1626908933
transform 1 0 29952 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_175
timestamp 1626908933
transform 1 0 30048 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_543
timestamp 1626908933
transform 1 0 30048 0 1 5328
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_161
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_431
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_161
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_431
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_161
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_431
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_171
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_459
timestamp 1626908933
transform 1 0 30600 0 1 5328
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_120
timestamp 1626908933
transform 1 0 30336 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_690
timestamp 1626908933
transform 1 0 30336 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_542
timestamp 1626908933
transform 1 0 31104 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_174
timestamp 1626908933
transform 1 0 31104 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_673
timestamp 1626908933
transform 1 0 31296 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_104
timestamp 1626908933
transform 1 0 31296 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_665
timestamp 1626908933
transform 1 0 31680 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_95
timestamp 1626908933
transform 1 0 31680 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_641
timestamp 1626908933
transform 1 0 32544 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_72
timestamp 1626908933
transform 1 0 32544 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_901
timestamp 1626908933
transform 1 0 32448 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_271
timestamp 1626908933
transform 1 0 32448 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_636
timestamp 1626908933
transform 1 0 32928 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_66
timestamp 1626908933
transform 1 0 32928 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_900
timestamp 1626908933
transform 1 0 33696 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_270
timestamp 1626908933
transform 1 0 33696 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_608
timestamp 1626908933
transform 1 0 33792 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_39
timestamp 1626908933
transform 1 0 33792 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_606
timestamp 1626908933
transform 1 0 34176 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_36
timestamp 1626908933
transform 1 0 34176 0 1 5328
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_416
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_146
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_416
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_146
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_416
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_146
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_155
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_443
timestamp 1626908933
transform 1 0 34600 0 1 5328
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_184
timestamp 1626908933
transform 1 0 34944 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_443
timestamp 1626908933
transform 1 0 34944 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_268
timestamp 1626908933
transform 1 0 35424 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_636
timestamp 1626908933
transform 1 0 35424 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_477
timestamp 1626908933
transform 1 0 35616 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1107
timestamp 1626908933
transform 1 0 35616 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_11
timestamp 1626908933
transform 1 0 35040 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_580
timestamp 1626908933
transform 1 0 35040 0 1 5328
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1483
timestamp 1626908933
transform 1 0 48 0 1 6179
box -32 -32 32 32
use M1M2_PR  M1M2_PR_715
timestamp 1626908933
transform 1 0 48 0 1 6179
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1530
timestamp 1626908933
transform 1 0 144 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_762
timestamp 1626908933
transform 1 0 144 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1108
timestamp 1626908933
transform 1 0 288 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_478
timestamp 1626908933
transform 1 0 288 0 -1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1572
timestamp 1626908933
transform 1 0 432 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_784
timestamp 1626908933
transform 1 0 432 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1199
timestamp 1626908933
transform 1 0 720 0 1 5883
box -29 -23 29 23
use L1M1_PR  L1M1_PR_411
timestamp 1626908933
transform 1 0 720 0 1 5883
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_400
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_130
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_400
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_130
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_400
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_130
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_427
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_139
timestamp 1626908933
transform 1 0 600 0 1 5994
box -200 -142 200 178
use L1M1_PR  L1M1_PR_782
timestamp 1626908933
transform 1 0 432 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1570
timestamp 1626908933
transform 1 0 432 0 1 6327
box -29 -23 29 23
use M1M2_PR  M1M2_PR_758
timestamp 1626908933
transform 1 0 336 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1526
timestamp 1626908933
transform 1 0 336 0 1 6327
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_24
timestamp 1626908933
transform 1 0 384 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_4
timestamp 1626908933
transform 1 0 384 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_559
timestamp 1626908933
transform 1 0 864 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1128
timestamp 1626908933
transform 1 0 864 0 -1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1099
timestamp 1626908933
transform 1 0 1200 0 1 5883
box -32 -32 32 32
use M1M2_PR  M1M2_PR_331
timestamp 1626908933
transform 1 0 1200 0 1 5883
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_541
timestamp 1626908933
transform 1 0 1248 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_173
timestamp 1626908933
transform 1 0 1248 0 -1 6660
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1067
timestamp 1626908933
transform 1 0 2064 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_299
timestamp 1626908933
transform 1 0 2064 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1069
timestamp 1626908933
transform 1 0 1584 0 1 5661
box -32 -32 32 32
use M1M2_PR  M1M2_PR_301
timestamp 1626908933
transform 1 0 1584 0 1 5661
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1132
timestamp 1626908933
transform 1 0 1440 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_562
timestamp 1626908933
transform 1 0 1440 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_540
timestamp 1626908933
transform 1 0 2208 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_172
timestamp 1626908933
transform 1 0 2208 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1109
timestamp 1626908933
transform 1 0 2400 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_479
timestamp 1626908933
transform 1 0 2400 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_442
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_183
timestamp 1626908933
transform 1 0 2496 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_539
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_171
timestamp 1626908933
transform 1 0 2592 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1114
timestamp 1626908933
transform 1 0 2784 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_545
timestamp 1626908933
transform 1 0 2784 0 -1 6660
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1156
timestamp 1626908933
transform 1 0 3120 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_368
timestamp 1626908933
transform 1 0 3120 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_942
timestamp 1626908933
transform 1 0 3312 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_154
timestamp 1626908933
transform 1 0 3312 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_890
timestamp 1626908933
transform 1 0 3504 0 1 5735
box -32 -32 32 32
use M1M2_PR  M1M2_PR_122
timestamp 1626908933
transform 1 0 3504 0 1 5735
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1155
timestamp 1626908933
transform 1 0 3600 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_367
timestamp 1626908933
transform 1 0 3600 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_936
timestamp 1626908933
transform 1 0 3792 0 1 5661
box -29 -23 29 23
use L1M1_PR  L1M1_PR_148
timestamp 1626908933
transform 1 0 3792 0 1 5661
box -29 -23 29 23
use M1M2_PR  M1M2_PR_121
timestamp 1626908933
transform 1 0 3504 0 1 6327
box -32 -32 32 32
use M1M2_PR  M1M2_PR_889
timestamp 1626908933
transform 1 0 3504 0 1 6327
box -32 -32 32 32
use L1M1_PR  L1M1_PR_149
timestamp 1626908933
transform 1 0 3504 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_365
timestamp 1626908933
transform 1 0 3312 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_937
timestamp 1626908933
transform 1 0 3504 0 1 6327
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1153
timestamp 1626908933
transform 1 0 3312 0 1 6327
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_99
timestamp 1626908933
transform 1 0 3168 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_44
timestamp 1626908933
transform 1 0 3168 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_526
timestamp 1626908933
transform 1 0 3648 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1095
timestamp 1626908933
transform 1 0 3648 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1107
timestamp 1626908933
transform 1 0 4032 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_537
timestamp 1626908933
transform 1 0 4032 0 -1 6660
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_385
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_115
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_385
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_115
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_385
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_115
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_123
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_411
timestamp 1626908933
transform 1 0 4600 0 1 5994
box -200 -142 200 178
use M1M2_PR  M1M2_PR_1479
timestamp 1626908933
transform 1 0 4272 0 1 6179
box -32 -32 32 32
use M1M2_PR  M1M2_PR_711
timestamp 1626908933
transform 1 0 4272 0 1 6179
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_269
timestamp 1626908933
transform 1 0 4800 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_899
timestamp 1626908933
transform 1 0 4800 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_518
timestamp 1626908933
transform 1 0 4896 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1087
timestamp 1626908933
transform 1 0 4896 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1093
timestamp 1626908933
transform 1 0 5280 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_523
timestamp 1626908933
transform 1 0 5280 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_898
timestamp 1626908933
transform 1 0 6048 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_268
timestamp 1626908933
transform 1 0 6048 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1067
timestamp 1626908933
transform 1 0 6144 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_498
timestamp 1626908933
transform 1 0 6144 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_897
timestamp 1626908933
transform 1 0 6528 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_267
timestamp 1626908933
transform 1 0 6528 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1079
timestamp 1626908933
transform 1 0 6624 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_509
timestamp 1626908933
transform 1 0 6624 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_895
timestamp 1626908933
transform 1 0 7776 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_265
timestamp 1626908933
transform 1 0 7776 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_896
timestamp 1626908933
transform 1 0 7392 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_266
timestamp 1626908933
transform 1 0 7392 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_538
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_170
timestamp 1626908933
transform 1 0 7584 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_441
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_182
timestamp 1626908933
transform 1 0 7488 0 -1 6660
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_100
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_370
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_100
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_370
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_100
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_370
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_107
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_395
timestamp 1626908933
transform 1 0 8600 0 1 5994
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_491
timestamp 1626908933
transform 1 0 7872 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1061
timestamp 1626908933
transform 1 0 7872 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1040
timestamp 1626908933
transform 1 0 8736 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_471
timestamp 1626908933
transform 1 0 8736 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1047
timestamp 1626908933
transform 1 0 9120 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_477
timestamp 1626908933
transform 1 0 9120 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_894
timestamp 1626908933
transform 1 0 8640 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_264
timestamp 1626908933
transform 1 0 8640 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1024
timestamp 1626908933
transform 1 0 9888 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_455
timestamp 1626908933
transform 1 0 9888 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_537
timestamp 1626908933
transform 1 0 10272 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_169
timestamp 1626908933
transform 1 0 10272 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1034
timestamp 1626908933
transform 1 0 10464 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_464
timestamp 1626908933
transform 1 0 10464 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_893
timestamp 1626908933
transform 1 0 11232 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_263
timestamp 1626908933
transform 1 0 11232 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_995
timestamp 1626908933
transform 1 0 11328 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_426
timestamp 1626908933
transform 1 0 11328 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1013
timestamp 1626908933
transform 1 0 11712 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_443
timestamp 1626908933
transform 1 0 11712 0 -1 6660
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_379
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_91
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_355
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_85
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_355
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_85
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_355
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_85
timestamp 1626908933
transform 1 0 12600 0 1 5994
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_968
timestamp 1626908933
transform 1 0 12576 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_399
timestamp 1626908933
transform 1 0 12576 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_440
timestamp 1626908933
transform 1 0 12480 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_181
timestamp 1626908933
transform 1 0 12480 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1000
timestamp 1626908933
transform 1 0 12960 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_430
timestamp 1626908933
transform 1 0 12960 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_947
timestamp 1626908933
transform 1 0 13920 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_378
timestamp 1626908933
transform 1 0 13920 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_536
timestamp 1626908933
transform 1 0 13728 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_168
timestamp 1626908933
transform 1 0 13728 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_986
timestamp 1626908933
transform 1 0 14304 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_416
timestamp 1626908933
transform 1 0 14304 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_892
timestamp 1626908933
transform 1 0 15072 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_262
timestamp 1626908933
transform 1 0 15072 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_928
timestamp 1626908933
transform 1 0 15168 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_359
timestamp 1626908933
transform 1 0 15168 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_966
timestamp 1626908933
transform 1 0 15552 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_396
timestamp 1626908933
transform 1 0 15552 0 -1 6660
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_70
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_340
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_70
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_340
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_70
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_340
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_75
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_363
timestamp 1626908933
transform 1 0 16600 0 1 5994
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_334
timestamp 1626908933
transform 1 0 16320 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_903
timestamp 1626908933
transform 1 0 16320 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_370
timestamp 1626908933
transform 1 0 16704 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_940
timestamp 1626908933
transform 1 0 16704 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_439
timestamp 1626908933
transform 1 0 17472 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_180
timestamp 1626908933
transform 1 0 17472 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_535
timestamp 1626908933
transform 1 0 17568 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_167
timestamp 1626908933
transform 1 0 17568 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_878
timestamp 1626908933
transform 1 0 17760 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_309
timestamp 1626908933
transform 1 0 17760 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_917
timestamp 1626908933
transform 1 0 18144 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_347
timestamp 1626908933
transform 1 0 18144 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_857
timestamp 1626908933
transform 1 0 18912 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_288
timestamp 1626908933
transform 1 0 18912 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_891
timestamp 1626908933
transform 1 0 19296 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_261
timestamp 1626908933
transform 1 0 19296 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_895
timestamp 1626908933
transform 1 0 19392 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_325
timestamp 1626908933
transform 1 0 19392 0 -1 6660
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_325
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_55
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_325
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_55
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_325
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_55
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_59
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_347
timestamp 1626908933
transform 1 0 20600 0 1 5994
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_534
timestamp 1626908933
transform 1 0 20160 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_166
timestamp 1626908933
transform 1 0 20160 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_272
timestamp 1626908933
transform 1 0 20352 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_841
timestamp 1626908933
transform 1 0 20352 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_863
timestamp 1626908933
transform 1 0 20736 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_293
timestamp 1626908933
transform 1 0 20736 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_533
timestamp 1626908933
transform 1 0 21504 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_165
timestamp 1626908933
transform 1 0 21504 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_839
timestamp 1626908933
transform 1 0 21696 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_269
timestamp 1626908933
transform 1 0 21696 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_890
timestamp 1626908933
transform 1 0 22560 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_260
timestamp 1626908933
transform 1 0 22560 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_825
timestamp 1626908933
transform 1 0 22656 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_255
timestamp 1626908933
transform 1 0 22656 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_438
timestamp 1626908933
transform 1 0 22464 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_179
timestamp 1626908933
transform 1 0 22464 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_790
timestamp 1626908933
transform 1 0 23424 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_221
timestamp 1626908933
transform 1 0 23424 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_889
timestamp 1626908933
transform 1 0 23808 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_259
timestamp 1626908933
transform 1 0 23808 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_802
timestamp 1626908933
transform 1 0 23904 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_232
timestamp 1626908933
transform 1 0 23904 0 -1 6660
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_331
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_43
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_310
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_40
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_310
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_40
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_310
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_40
timestamp 1626908933
transform 1 0 24600 0 1 5994
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_532
timestamp 1626908933
transform 1 0 24672 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_164
timestamp 1626908933
transform 1 0 24672 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_202
timestamp 1626908933
transform 1 0 24864 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_771
timestamp 1626908933
transform 1 0 24864 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_781
timestamp 1626908933
transform 1 0 25248 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_211
timestamp 1626908933
transform 1 0 25248 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_753
timestamp 1626908933
transform 1 0 26016 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_184
timestamp 1626908933
transform 1 0 26016 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_888
timestamp 1626908933
transform 1 0 26400 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_258
timestamp 1626908933
transform 1 0 26400 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_759
timestamp 1626908933
transform 1 0 26496 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_189
timestamp 1626908933
transform 1 0 26496 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_163
timestamp 1626908933
transform 1 0 27552 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_531
timestamp 1626908933
transform 1 0 27552 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_178
timestamp 1626908933
transform 1 0 27456 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_437
timestamp 1626908933
transform 1 0 27456 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_257
timestamp 1626908933
transform 1 0 27264 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_480
timestamp 1626908933
transform 1 0 27360 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_887
timestamp 1626908933
transform 1 0 27264 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1110
timestamp 1626908933
transform 1 0 27360 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_256
timestamp 1626908933
transform 1 0 27744 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_886
timestamp 1626908933
transform 1 0 27744 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_167
timestamp 1626908933
transform 1 0 27840 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_737
timestamp 1626908933
transform 1 0 27840 0 -1 6660
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_315
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_27
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_25
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_295
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_25
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_295
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_25
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_295
timestamp 1626908933
transform 1 0 28600 0 1 5994
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_147
timestamp 1626908933
transform 1 0 28608 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_716
timestamp 1626908933
transform 1 0 28608 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_885
timestamp 1626908933
transform 1 0 28992 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_255
timestamp 1626908933
transform 1 0 28992 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_713
timestamp 1626908933
transform 1 0 29088 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_143
timestamp 1626908933
transform 1 0 29088 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_884
timestamp 1626908933
transform 1 0 29856 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_254
timestamp 1626908933
transform 1 0 29856 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_691
timestamp 1626908933
transform 1 0 29952 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_122
timestamp 1626908933
transform 1 0 29952 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_689
timestamp 1626908933
transform 1 0 30336 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_119
timestamp 1626908933
transform 1 0 30336 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_530
timestamp 1626908933
transform 1 0 31104 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_162
timestamp 1626908933
transform 1 0 31104 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_672
timestamp 1626908933
transform 1 0 31296 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_103
timestamp 1626908933
transform 1 0 31296 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_664
timestamp 1626908933
transform 1 0 31680 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_94
timestamp 1626908933
transform 1 0 31680 0 -1 6660
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_299
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_11
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_280
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_10
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_280
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_10
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_280
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_10
timestamp 1626908933
transform 1 0 32600 0 1 5994
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_436
timestamp 1626908933
transform 1 0 32448 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_177
timestamp 1626908933
transform 1 0 32448 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_71
timestamp 1626908933
transform 1 0 32544 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_640
timestamp 1626908933
transform 1 0 32544 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_635
timestamp 1626908933
transform 1 0 32928 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_65
timestamp 1626908933
transform 1 0 32928 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_883
timestamp 1626908933
transform 1 0 33696 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_253
timestamp 1626908933
transform 1 0 33696 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_607
timestamp 1626908933
transform 1 0 33792 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_38
timestamp 1626908933
transform 1 0 33792 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_605
timestamp 1626908933
transform 1 0 34176 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_35
timestamp 1626908933
transform 1 0 34176 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_10
timestamp 1626908933
transform 1 0 34944 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_580
timestamp 1626908933
transform 1 0 34944 0 -1 6660
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1436
timestamp 1626908933
transform 1 0 144 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_668
timestamp 1626908933
transform 1 0 144 0 1 6919
box -32 -32 32 32
use M2M3_PR  M2M3_PR_113
timestamp 1626908933
transform 1 0 48 0 1 6503
box -33 -37 33 37
use M2M3_PR  M2M3_PR_54
timestamp 1626908933
transform 1 0 48 0 1 6503
box -33 -37 33 37
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_435
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_176
timestamp 1626908933
transform 1 0 288 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_481
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1111
timestamp 1626908933
transform 1 0 384 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_402
timestamp 1626908933
transform 1 0 336 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1170
timestamp 1626908933
transform 1 0 336 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_700
timestamp 1626908933
transform 1 0 528 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1488
timestamp 1626908933
transform 1 0 528 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_369
timestamp 1626908933
transform 1 0 720 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_423
timestamp 1626908933
transform 1 0 720 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1157
timestamp 1626908933
transform 1 0 720 0 1 6771
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1211
timestamp 1626908933
transform 1 0 720 0 1 6549
box -29 -23 29 23
use L1M1_PR  L1M1_PR_409
timestamp 1626908933
transform 1 0 816 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_470
timestamp 1626908933
transform 1 0 624 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1197
timestamp 1626908933
transform 1 0 816 0 1 6919
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1258
timestamp 1626908933
transform 1 0 624 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_558
timestamp 1626908933
transform 1 0 864 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1127
timestamp 1626908933
transform 1 0 864 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_1
timestamp 1626908933
transform 1 0 480 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_26
timestamp 1626908933
transform 1 0 480 0 1 6660
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1098
timestamp 1626908933
transform 1 0 1200 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_330
timestamp 1626908933
transform 1 0 1200 0 1 6919
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1117
timestamp 1626908933
transform 1 0 1392 0 1 6549
box -32 -32 32 32
use M1M2_PR  M1M2_PR_349
timestamp 1626908933
transform 1 0 1392 0 1 6549
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_5
timestamp 1626908933
transform 1 0 1248 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_25
timestamp 1626908933
transform 1 0 1248 0 1 6660
box -38 -49 518 715
use M1M2_PR  M1M2_PR_300
timestamp 1626908933
transform 1 0 1584 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1068
timestamp 1626908933
transform 1 0 1584 0 1 6771
box -32 -32 32 32
use M1M2_PR  M1M2_PR_764
timestamp 1626908933
transform 1 0 1776 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1532
timestamp 1626908933
transform 1 0 1776 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_786
timestamp 1626908933
transform 1 0 1584 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1574
timestamp 1626908933
transform 1 0 1584 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_556
timestamp 1626908933
transform 1 0 2112 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1126
timestamp 1626908933
transform 1 0 2112 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_551
timestamp 1626908933
transform 1 0 1728 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1120
timestamp 1626908933
transform 1 0 1728 0 1 6660
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_570
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_282
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_265
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_535
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_265
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_535
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_265
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_535
timestamp 1626908933
transform 1 0 2600 0 1 6660
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_482
timestamp 1626908933
transform 1 0 2880 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1112
timestamp 1626908933
transform 1 0 2880 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_102
timestamp 1626908933
transform 1 0 2976 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_47
timestamp 1626908933
transform 1 0 2976 0 1 6660
box -38 -49 518 715
use L1M1_PR  L1M1_PR_373
timestamp 1626908933
transform 1 0 3216 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1161
timestamp 1626908933
transform 1 0 3216 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_120
timestamp 1626908933
transform 1 0 3504 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_888
timestamp 1626908933
transform 1 0 3504 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_153
timestamp 1626908933
transform 1 0 3312 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_941
timestamp 1626908933
transform 1 0 3312 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_252
timestamp 1626908933
transform 1 0 3936 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_882
timestamp 1626908933
transform 1 0 3936 0 1 6660
box -38 -49 134 715
use L1M1_PR  L1M1_PR_147
timestamp 1626908933
transform 1 0 3792 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_935
timestamp 1626908933
transform 1 0 3792 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_302
timestamp 1626908933
transform 1 0 3600 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1070
timestamp 1626908933
transform 1 0 3600 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_370
timestamp 1626908933
transform 1 0 3600 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1158
timestamp 1626908933
transform 1 0 3600 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_103
timestamp 1626908933
transform 1 0 3456 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_48
timestamp 1626908933
transform 1 0 3456 0 1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1106
timestamp 1626908933
transform 1 0 4032 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_536
timestamp 1626908933
transform 1 0 4032 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_529
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_161
timestamp 1626908933
transform 1 0 5088 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1113
timestamp 1626908933
transform 1 0 4896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_881
timestamp 1626908933
transform 1 0 4800 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_483
timestamp 1626908933
transform 1 0 4896 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_251
timestamp 1626908933
transform 1 0 4800 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_434
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_175
timestamp 1626908933
transform 1 0 4992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_515
timestamp 1626908933
transform 1 0 5376 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1084
timestamp 1626908933
transform 1 0 5376 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_250
timestamp 1626908933
transform 1 0 5280 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_880
timestamp 1626908933
transform 1 0 5280 0 1 6660
box -38 -49 134 715
use M1M2_PR  M1M2_PR_747
timestamp 1626908933
transform 1 0 5424 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1515
timestamp 1626908933
transform 1 0 5424 0 1 6993
box -32 -32 32 32
use L1M1_PR  L1M1_PR_773
timestamp 1626908933
transform 1 0 5904 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1561
timestamp 1626908933
transform 1 0 5904 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_76
timestamp 1626908933
transform 1 0 5760 0 1 6660
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_156
timestamp 1626908933
transform 1 0 5760 0 1 6660
box -38 -49 902 715
use osc_core_VIA4  osc_core_VIA4_554
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_266
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_250
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_520
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_250
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_520
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_250
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_520
timestamp 1626908933
transform 1 0 6600 0 1 6660
box -200 -49 200 49
use L1M1_PR  L1M1_PR_140
timestamp 1626908933
transform 1 0 6288 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_928
timestamp 1626908933
transform 1 0 6288 0 1 6993
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_508
timestamp 1626908933
transform 1 0 6624 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1078
timestamp 1626908933
transform 1 0 6624 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_879
timestamp 1626908933
transform 1 0 7392 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_249
timestamp 1626908933
transform 1 0 7392 0 1 6660
box -38 -49 134 715
use M2M3_PR  M2M3_PR_112
timestamp 1626908933
transform 1 0 7632 0 1 6503
box -33 -37 33 37
use M2M3_PR  M2M3_PR_53
timestamp 1626908933
transform 1 0 7632 0 1 6503
box -33 -37 33 37
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1055
timestamp 1626908933
transform 1 0 7488 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_486
timestamp 1626908933
transform 1 0 7488 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1060
timestamp 1626908933
transform 1 0 7872 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_490
timestamp 1626908933
transform 1 0 7872 0 1 6660
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1522
timestamp 1626908933
transform 1 0 8784 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_734
timestamp 1626908933
transform 1 0 8784 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1476
timestamp 1626908933
transform 1 0 7920 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_708
timestamp 1626908933
transform 1 0 7920 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_149
timestamp 1626908933
transform 1 0 8640 0 1 6660
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_69
timestamp 1626908933
transform 1 0 8640 0 1 6660
box -38 -49 902 715
use L1M1_PR  L1M1_PR_913
timestamp 1626908933
transform 1 0 9168 0 1 6993
box -29 -23 29 23
use L1M1_PR  L1M1_PR_125
timestamp 1626908933
transform 1 0 9168 0 1 6993
box -29 -23 29 23
use M1M2_PR  M1M2_PR_875
timestamp 1626908933
transform 1 0 9168 0 1 6993
box -32 -32 32 32
use M1M2_PR  M1M2_PR_107
timestamp 1626908933
transform 1 0 9168 0 1 6993
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1036
timestamp 1626908933
transform 1 0 9504 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_467
timestamp 1626908933
transform 1 0 9504 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_174
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_433
timestamp 1626908933
transform 1 0 9984 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_484
timestamp 1626908933
transform 1 0 9888 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1114
timestamp 1626908933
transform 1 0 9888 0 1 6660
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_538
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_250
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_235
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_505
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_235
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_505
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_235
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_505
timestamp 1626908933
transform 1 0 10600 0 1 6660
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_463
timestamp 1626908933
transform 1 0 10464 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1033
timestamp 1626908933
transform 1 0 10464 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_448
timestamp 1626908933
transform 1 0 10080 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1017
timestamp 1626908933
transform 1 0 10080 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_878
timestamp 1626908933
transform 1 0 11232 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_248
timestamp 1626908933
transform 1 0 11232 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_994
timestamp 1626908933
transform 1 0 11328 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_425
timestamp 1626908933
transform 1 0 11328 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1012
timestamp 1626908933
transform 1 0 11712 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_442
timestamp 1626908933
transform 1 0 11712 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_976
timestamp 1626908933
transform 1 0 12480 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_407
timestamp 1626908933
transform 1 0 12480 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_877
timestamp 1626908933
transform 1 0 12864 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_247
timestamp 1626908933
transform 1 0 12864 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_999
timestamp 1626908933
transform 1 0 12960 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_429
timestamp 1626908933
transform 1 0 12960 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_876
timestamp 1626908933
transform 1 0 13728 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_246
timestamp 1626908933
transform 1 0 13728 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_946
timestamp 1626908933
transform 1 0 13824 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_377
timestamp 1626908933
transform 1 0 13824 0 1 6660
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_522
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_234
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_220
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_490
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_220
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_490
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_220
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_490
timestamp 1626908933
transform 1 0 14600 0 1 6660
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_173
timestamp 1626908933
transform 1 0 14976 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_432
timestamp 1626908933
transform 1 0 14976 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_415
timestamp 1626908933
transform 1 0 14208 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_985
timestamp 1626908933
transform 1 0 14208 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_875
timestamp 1626908933
transform 1 0 15072 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_245
timestamp 1626908933
transform 1 0 15072 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_927
timestamp 1626908933
transform 1 0 15168 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_358
timestamp 1626908933
transform 1 0 15168 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_965
timestamp 1626908933
transform 1 0 15552 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_395
timestamp 1626908933
transform 1 0 15552 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_939
timestamp 1626908933
transform 1 0 16896 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_369
timestamp 1626908933
transform 1 0 16896 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_528
timestamp 1626908933
transform 1 0 16320 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_160
timestamp 1626908933
transform 1 0 16320 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_902
timestamp 1626908933
transform 1 0 16512 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_333
timestamp 1626908933
transform 1 0 16512 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_874
timestamp 1626908933
transform 1 0 17664 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_244
timestamp 1626908933
transform 1 0 17664 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_877
timestamp 1626908933
transform 1 0 17760 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_308
timestamp 1626908933
transform 1 0 17760 0 1 6660
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_506
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_218
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_205
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_475
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_205
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_475
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_205
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_475
timestamp 1626908933
transform 1 0 18600 0 1 6660
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_346
timestamp 1626908933
transform 1 0 18144 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_916
timestamp 1626908933
transform 1 0 18144 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_873
timestamp 1626908933
transform 1 0 19104 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_243
timestamp 1626908933
transform 1 0 19104 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_527
timestamp 1626908933
transform 1 0 18912 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_159
timestamp 1626908933
transform 1 0 18912 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_894
timestamp 1626908933
transform 1 0 19200 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_324
timestamp 1626908933
transform 1 0 19200 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_874
timestamp 1626908933
transform 1 0 20064 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_304
timestamp 1626908933
transform 1 0 20064 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_431
timestamp 1626908933
transform 1 0 19968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_172
timestamp 1626908933
transform 1 0 19968 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_526
timestamp 1626908933
transform 1 0 20832 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_158
timestamp 1626908933
transform 1 0 20832 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_825
timestamp 1626908933
transform 1 0 21024 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_256
timestamp 1626908933
transform 1 0 21024 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_848
timestamp 1626908933
transform 1 0 21408 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_278
timestamp 1626908933
transform 1 0 21408 0 1 6660
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_490
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_202
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_460
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_190
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_460
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_190
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_460
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_190
timestamp 1626908933
transform 1 0 22600 0 1 6660
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_872
timestamp 1626908933
transform 1 0 22176 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_242
timestamp 1626908933
transform 1 0 22176 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_237
timestamp 1626908933
transform 1 0 22272 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_806
timestamp 1626908933
transform 1 0 22272 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_824
timestamp 1626908933
transform 1 0 22656 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_254
timestamp 1626908933
transform 1 0 22656 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_789
timestamp 1626908933
transform 1 0 23424 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_220
timestamp 1626908933
transform 1 0 23424 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_871
timestamp 1626908933
transform 1 0 23808 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_241
timestamp 1626908933
transform 1 0 23808 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_801
timestamp 1626908933
transform 1 0 23904 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_231
timestamp 1626908933
transform 1 0 23904 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_525
timestamp 1626908933
transform 1 0 25056 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_157
timestamp 1626908933
transform 1 0 25056 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_430
timestamp 1626908933
transform 1 0 24960 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_171
timestamp 1626908933
transform 1 0 24960 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_637
timestamp 1626908933
transform 1 0 24672 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_269
timestamp 1626908933
transform 1 0 24672 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1115
timestamp 1626908933
transform 1 0 24864 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_485
timestamp 1626908933
transform 1 0 24864 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_780
timestamp 1626908933
transform 1 0 25248 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_210
timestamp 1626908933
transform 1 0 25248 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_752
timestamp 1626908933
transform 1 0 26016 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_183
timestamp 1626908933
transform 1 0 26016 0 1 6660
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_474
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_186
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_445
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_175
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_445
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_175
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_445
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_175
timestamp 1626908933
transform 1 0 26600 0 1 6660
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_870
timestamp 1626908933
transform 1 0 26400 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_240
timestamp 1626908933
transform 1 0 26400 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_188
timestamp 1626908933
transform 1 0 26496 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_758
timestamp 1626908933
transform 1 0 26496 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_736
timestamp 1626908933
transform 1 0 27840 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_166
timestamp 1626908933
transform 1 0 27840 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_524
timestamp 1626908933
transform 1 0 27264 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_156
timestamp 1626908933
transform 1 0 27264 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_733
timestamp 1626908933
transform 1 0 27456 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_164
timestamp 1626908933
transform 1 0 27456 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_715
timestamp 1626908933
transform 1 0 28608 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_146
timestamp 1626908933
transform 1 0 28608 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_869
timestamp 1626908933
transform 1 0 28992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_239
timestamp 1626908933
transform 1 0 28992 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_712
timestamp 1626908933
transform 1 0 29088 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_142
timestamp 1626908933
transform 1 0 29088 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1116
timestamp 1626908933
transform 1 0 29856 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_486
timestamp 1626908933
transform 1 0 29856 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_238
timestamp 1626908933
transform 1 0 30240 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_868
timestamp 1626908933
transform 1 0 30240 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_170
timestamp 1626908933
transform 1 0 29952 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_429
timestamp 1626908933
transform 1 0 29952 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_155
timestamp 1626908933
transform 1 0 30048 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_523
timestamp 1626908933
transform 1 0 30048 0 1 6660
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_160
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_430
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_160
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_430
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_160
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_430
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_170
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_458
timestamp 1626908933
transform 1 0 30600 0 1 6660
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_118
timestamp 1626908933
transform 1 0 30336 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_688
timestamp 1626908933
transform 1 0 30336 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_522
timestamp 1626908933
transform 1 0 31104 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_154
timestamp 1626908933
transform 1 0 31104 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_671
timestamp 1626908933
transform 1 0 31296 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_102
timestamp 1626908933
transform 1 0 31296 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_663
timestamp 1626908933
transform 1 0 31680 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_93
timestamp 1626908933
transform 1 0 31680 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_867
timestamp 1626908933
transform 1 0 32448 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_237
timestamp 1626908933
transform 1 0 32448 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_639
timestamp 1626908933
transform 1 0 32544 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_70
timestamp 1626908933
transform 1 0 32544 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_634
timestamp 1626908933
transform 1 0 32928 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_64
timestamp 1626908933
transform 1 0 32928 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_866
timestamp 1626908933
transform 1 0 33696 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_236
timestamp 1626908933
transform 1 0 33696 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_606
timestamp 1626908933
transform 1 0 33792 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_37
timestamp 1626908933
transform 1 0 33792 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_604
timestamp 1626908933
transform 1 0 34176 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_34
timestamp 1626908933
transform 1 0 34176 0 1 6660
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_415
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_145
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_415
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_145
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_415
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_145
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_154
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_442
timestamp 1626908933
transform 1 0 34600 0 1 6660
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_169
timestamp 1626908933
transform 1 0 34944 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_428
timestamp 1626908933
transform 1 0 34944 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_10
timestamp 1626908933
transform 1 0 35040 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_579
timestamp 1626908933
transform 1 0 35040 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_270
timestamp 1626908933
transform 1 0 35424 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_638
timestamp 1626908933
transform 1 0 35424 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_487
timestamp 1626908933
transform 1 0 35616 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1117
timestamp 1626908933
transform 1 0 35616 0 1 6660
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_399
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_129
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_399
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_129
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_399
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_129
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1489
timestamp 1626908933
transform 1 0 432 0 1 7437
box -29 -23 29 23
use L1M1_PR  L1M1_PR_701
timestamp 1626908933
transform 1 0 432 0 1 7437
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1437
timestamp 1626908933
transform 1 0 240 0 1 7437
box -32 -32 32 32
use M1M2_PR  M1M2_PR_669
timestamp 1626908933
transform 1 0 240 0 1 7437
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_426
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_138
timestamp 1626908933
transform 1 0 600 0 1 7326
box -200 -142 200 178
use M1M2_PR  M1M2_PR_401
timestamp 1626908933
transform 1 0 336 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1169
timestamp 1626908933
transform 1 0 336 0 1 7659
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_271
timestamp 1626908933
transform 1 0 288 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_639
timestamp 1626908933
transform 1 0 288 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_2
timestamp 1626908933
transform 1 0 480 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_27
timestamp 1626908933
transform 1 0 480 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1257
timestamp 1626908933
transform 1 0 624 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1204
timestamp 1626908933
transform 1 0 816 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_469
timestamp 1626908933
transform 1 0 624 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_416
timestamp 1626908933
transform 1 0 816 0 1 7733
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1126
timestamp 1626908933
transform 1 0 864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_557
timestamp 1626908933
transform 1 0 864 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1162
timestamp 1626908933
transform 1 0 816 0 1 7585
box -29 -23 29 23
use L1M1_PR  L1M1_PR_374
timestamp 1626908933
transform 1 0 816 0 1 7585
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1109
timestamp 1626908933
transform 1 0 1008 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_341
timestamp 1626908933
transform 1 0 1008 0 1 7733
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_521
timestamp 1626908933
transform 1 0 1248 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_153
timestamp 1626908933
transform 1 0 1248 0 -1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_357
timestamp 1626908933
transform 1 0 1776 0 1 7215
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1125
timestamp 1626908933
transform 1 0 1776 0 1 7215
box -32 -32 32 32
use L1M1_PR  L1M1_PR_429
timestamp 1626908933
transform 1 0 1584 0 1 7215
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1217
timestamp 1626908933
transform 1 0 1584 0 1 7215
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_152
timestamp 1626908933
transform 1 0 2208 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_520
timestamp 1626908933
transform 1 0 2208 0 -1 7992
box -38 -49 230 715
use M1M2_PR  M1M2_PR_297
timestamp 1626908933
transform 1 0 2256 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1065
timestamp 1626908933
transform 1 0 2256 0 1 7733
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_561
timestamp 1626908933
transform 1 0 1440 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1131
timestamp 1626908933
transform 1 0 1440 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_168
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_427
timestamp 1626908933
transform 1 0 2496 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_488
timestamp 1626908933
transform 1 0 2400 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1118
timestamp 1626908933
transform 1 0 2400 0 -1 7992
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_569
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_281
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_4
timestamp 1626908933
transform 1 0 2976 0 -1 7992
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_9
timestamp 1626908933
transform 1 0 2976 0 -1 7992
box -38 -49 326 715
use L1M1_PR  L1M1_PR_363
timestamp 1626908933
transform 1 0 3024 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1151
timestamp 1626908933
transform 1 0 3024 0 1 7733
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_544
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1113
timestamp 1626908933
transform 1 0 2592 0 -1 7992
box -38 -49 422 715
use L1M1_PR  L1M1_PR_938
timestamp 1626908933
transform 1 0 3408 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_150
timestamp 1626908933
transform 1 0 3408 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1159
timestamp 1626908933
transform 1 0 3504 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_371
timestamp 1626908933
transform 1 0 3504 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1072
timestamp 1626908933
transform 1 0 3504 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_304
timestamp 1626908933
transform 1 0 3504 0 1 7659
box -32 -32 32 32
use L1M1_PR  L1M1_PR_943
timestamp 1626908933
transform 1 0 3216 0 1 7733
box -29 -23 29 23
use L1M1_PR  L1M1_PR_155
timestamp 1626908933
transform 1 0 3216 0 1 7733
box -29 -23 29 23
use M1M2_PR  M1M2_PR_894
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_126
timestamp 1626908933
transform 1 0 3312 0 1 7733
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_151
timestamp 1626908933
transform 1 0 3744 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_519
timestamp 1626908933
transform 1 0 3744 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_235
timestamp 1626908933
transform 1 0 3936 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_865
timestamp 1626908933
transform 1 0 3936 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_105
timestamp 1626908933
transform -1 0 3744 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_50
timestamp 1626908933
transform -1 0 3744 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1105
timestamp 1626908933
transform 1 0 4032 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_535
timestamp 1626908933
transform 1 0 4032 0 -1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_410
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_122
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_114
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_384
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_114
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_384
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_114
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_384
timestamp 1626908933
transform 1 0 4600 0 1 7326
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_150
timestamp 1626908933
transform 1 0 4800 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_518
timestamp 1626908933
transform 1 0 4800 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_522
timestamp 1626908933
transform 1 0 4992 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1092
timestamp 1626908933
transform 1 0 4992 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1560
timestamp 1626908933
transform 1 0 5904 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_772
timestamp 1626908933
transform 1 0 5904 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1514
timestamp 1626908933
transform 1 0 5424 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_746
timestamp 1626908933
transform 1 0 5424 0 1 7659
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_159
timestamp 1626908933
transform 1 0 5760 0 -1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_79
timestamp 1626908933
transform 1 0 5760 0 -1 7992
box -38 -49 902 715
use M1M2_PR  M1M2_PR_886
timestamp 1626908933
transform 1 0 6288 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_118
timestamp 1626908933
transform 1 0 6288 0 1 7659
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_265
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_553
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -142 200 178
use L1M1_PR  L1M1_PR_927
timestamp 1626908933
transform 1 0 6480 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_139
timestamp 1626908933
transform 1 0 6480 0 1 7659
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1077
timestamp 1626908933
transform 1 0 6624 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_507
timestamp 1626908933
transform 1 0 6624 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_489
timestamp 1626908933
transform 1 0 7392 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1119
timestamp 1626908933
transform 1 0 7392 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_167
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_426
timestamp 1626908933
transform 1 0 7488 0 -1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_737
timestamp 1626908933
transform 1 0 7824 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1525
timestamp 1626908933
transform 1 0 7824 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_689
timestamp 1626908933
transform 1 0 7632 0 1 7807
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1457
timestamp 1626908933
transform 1 0 7632 0 1 7807
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_70
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_150
timestamp 1626908933
transform 1 0 7584 0 -1 7992
box -38 -49 902 715
use M1M2_PR  M1M2_PR_1475
timestamp 1626908933
transform 1 0 7920 0 1 7733
box -32 -32 32 32
use M1M2_PR  M1M2_PR_707
timestamp 1626908933
transform 1 0 7920 0 1 7733
box -32 -32 32 32
use L1M1_PR  L1M1_PR_922
timestamp 1626908933
transform 1 0 8112 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_134
timestamp 1626908933
transform 1 0 8112 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_883
timestamp 1626908933
transform 1 0 8112 0 1 7659
box -32 -32 32 32
use M1M2_PR  M1M2_PR_115
timestamp 1626908933
transform 1 0 8112 0 1 7659
box -32 -32 32 32
use M3M4_PR  M3M4_PR_33
timestamp 1626908933
transform 1 0 8112 0 1 7601
box -38 -33 38 33
use M3M4_PR  M3M4_PR_12
timestamp 1626908933
transform 1 0 8112 0 1 7601
box -38 -33 38 33
use M2M3_PR  M2M3_PR_72
timestamp 1626908933
transform 1 0 8112 0 1 7601
box -33 -37 33 37
use M2M3_PR  M2M3_PR_13
timestamp 1626908933
transform 1 0 8112 0 1 7601
box -33 -37 33 37
use osc_core_VIA4  osc_core_VIA4_394
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_106
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_369
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_99
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_369
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_99
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_369
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_99
timestamp 1626908933
transform 1 0 8600 0 1 7326
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1120
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_490
timestamp 1626908933
transform 1 0 8640 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_640
timestamp 1626908933
transform 1 0 8448 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_272
timestamp 1626908933
transform 1 0 8448 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_66
timestamp 1626908933
transform 1 0 8736 0 -1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_146
timestamp 1626908933
transform 1 0 8736 0 -1 7992
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1507
timestamp 1626908933
transform 1 0 8880 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_912
timestamp 1626908933
transform 1 0 9264 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_719
timestamp 1626908933
transform 1 0 8880 0 1 7659
box -29 -23 29 23
use L1M1_PR  L1M1_PR_124
timestamp 1626908933
transform 1 0 9264 0 1 7659
box -29 -23 29 23
use M1M2_PR  M1M2_PR_874
timestamp 1626908933
transform 1 0 9168 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_106
timestamp 1626908933
transform 1 0 9168 0 1 7585
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_517
timestamp 1626908933
transform 1 0 9600 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_149
timestamp 1626908933
transform 1 0 9600 0 -1 7992
box -38 -49 230 715
use osc_core_VIA4  osc_core_VIA4_249
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_537
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1045
timestamp 1626908933
transform 1 0 9792 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_475
timestamp 1626908933
transform 1 0 9792 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_864
timestamp 1626908933
transform 1 0 10560 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_234
timestamp 1626908933
transform 1 0 10560 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1009
timestamp 1626908933
transform 1 0 10656 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_440
timestamp 1626908933
transform 1 0 10656 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1026
timestamp 1626908933
transform 1 0 11040 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_456
timestamp 1626908933
transform 1 0 11040 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_516
timestamp 1626908933
transform 1 0 11808 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_148
timestamp 1626908933
transform 1 0 11808 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_989
timestamp 1626908933
transform 1 0 12096 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_420
timestamp 1626908933
transform 1 0 12096 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_863
timestamp 1626908933
transform 1 0 12000 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_233
timestamp 1626908933
transform 1 0 12000 0 -1 7992
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_378
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_90
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_354
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_84
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_354
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_84
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_354
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_84
timestamp 1626908933
transform 1 0 12600 0 1 7326
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_967
timestamp 1626908933
transform 1 0 12576 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_398
timestamp 1626908933
transform 1 0 12576 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_425
timestamp 1626908933
transform 1 0 12480 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_166
timestamp 1626908933
transform 1 0 12480 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_998
timestamp 1626908933
transform 1 0 12960 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_428
timestamp 1626908933
transform 1 0 12960 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_945
timestamp 1626908933
transform 1 0 13920 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_376
timestamp 1626908933
transform 1 0 13920 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_515
timestamp 1626908933
transform 1 0 13728 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_147
timestamp 1626908933
transform 1 0 13728 0 -1 7992
box -38 -49 230 715
use osc_core_VIA4  osc_core_VIA4_233
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_521
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_984
timestamp 1626908933
transform 1 0 14304 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_414
timestamp 1626908933
transform 1 0 14304 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_862
timestamp 1626908933
transform 1 0 15072 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_232
timestamp 1626908933
transform 1 0 15072 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_926
timestamp 1626908933
transform 1 0 15168 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_357
timestamp 1626908933
transform 1 0 15168 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_964
timestamp 1626908933
transform 1 0 15552 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_394
timestamp 1626908933
transform 1 0 15552 0 -1 7992
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1348
timestamp 1626908933
transform 1 0 15792 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_580
timestamp 1626908933
transform 1 0 15792 0 1 7585
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_69
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_339
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_69
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_339
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_69
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_339
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_74
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_362
timestamp 1626908933
transform 1 0 16600 0 1 7326
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_332
timestamp 1626908933
transform 1 0 16320 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_901
timestamp 1626908933
transform 1 0 16320 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_368
timestamp 1626908933
transform 1 0 16704 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_938
timestamp 1626908933
transform 1 0 16704 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_424
timestamp 1626908933
transform 1 0 17472 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_165
timestamp 1626908933
transform 1 0 17472 0 -1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1346
timestamp 1626908933
transform 1 0 17616 0 1 7585
box -32 -32 32 32
use M1M2_PR  M1M2_PR_578
timestamp 1626908933
transform 1 0 17616 0 1 7585
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_514
timestamp 1626908933
transform 1 0 17568 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_146
timestamp 1626908933
transform 1 0 17568 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_876
timestamp 1626908933
transform 1 0 17760 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_307
timestamp 1626908933
transform 1 0 17760 0 -1 7992
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_217
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_505
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_915
timestamp 1626908933
transform 1 0 18144 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_345
timestamp 1626908933
transform 1 0 18144 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_856
timestamp 1626908933
transform 1 0 18912 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_287
timestamp 1626908933
transform 1 0 18912 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_861
timestamp 1626908933
transform 1 0 19296 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_231
timestamp 1626908933
transform 1 0 19296 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_893
timestamp 1626908933
transform 1 0 19392 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_323
timestamp 1626908933
transform 1 0 19392 0 -1 7992
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_324
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_54
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_324
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_54
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_324
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_54
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_58
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_346
timestamp 1626908933
transform 1 0 20600 0 1 7326
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_513
timestamp 1626908933
transform 1 0 20160 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_145
timestamp 1626908933
transform 1 0 20160 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_271
timestamp 1626908933
transform 1 0 20352 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_840
timestamp 1626908933
transform 1 0 20352 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_862
timestamp 1626908933
transform 1 0 20736 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_292
timestamp 1626908933
transform 1 0 20736 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_512
timestamp 1626908933
transform 1 0 21504 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_144
timestamp 1626908933
transform 1 0 21504 0 -1 7992
box -38 -49 230 715
use osc_core_VIA4  osc_core_VIA4_489
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_201
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_838
timestamp 1626908933
transform 1 0 21696 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_268
timestamp 1626908933
transform 1 0 21696 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_860
timestamp 1626908933
transform 1 0 22560 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_230
timestamp 1626908933
transform 1 0 22560 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_823
timestamp 1626908933
transform 1 0 22656 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_253
timestamp 1626908933
transform 1 0 22656 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_423
timestamp 1626908933
transform 1 0 22464 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_164
timestamp 1626908933
transform 1 0 22464 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_788
timestamp 1626908933
transform 1 0 23424 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_219
timestamp 1626908933
transform 1 0 23424 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_859
timestamp 1626908933
transform 1 0 23808 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_229
timestamp 1626908933
transform 1 0 23808 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_800
timestamp 1626908933
transform 1 0 23904 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_230
timestamp 1626908933
transform 1 0 23904 0 -1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_330
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_42
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_309
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_39
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_309
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_39
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_309
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_39
timestamp 1626908933
transform 1 0 24600 0 1 7326
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_511
timestamp 1626908933
transform 1 0 24672 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_143
timestamp 1626908933
transform 1 0 24672 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_201
timestamp 1626908933
transform 1 0 24864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_770
timestamp 1626908933
transform 1 0 24864 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_779
timestamp 1626908933
transform 1 0 25248 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_209
timestamp 1626908933
transform 1 0 25248 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_751
timestamp 1626908933
transform 1 0 26016 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_182
timestamp 1626908933
transform 1 0 26016 0 -1 7992
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_473
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_185
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_858
timestamp 1626908933
transform 1 0 26400 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_228
timestamp 1626908933
transform 1 0 26400 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_757
timestamp 1626908933
transform 1 0 26496 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_187
timestamp 1626908933
transform 1 0 26496 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_142
timestamp 1626908933
transform 1 0 27552 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_510
timestamp 1626908933
transform 1 0 27552 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_163
timestamp 1626908933
transform 1 0 27456 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_422
timestamp 1626908933
transform 1 0 27456 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_227
timestamp 1626908933
transform 1 0 27264 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_491
timestamp 1626908933
transform 1 0 27360 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_857
timestamp 1626908933
transform 1 0 27264 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1121
timestamp 1626908933
transform 1 0 27360 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_226
timestamp 1626908933
transform 1 0 27744 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_856
timestamp 1626908933
transform 1 0 27744 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_165
timestamp 1626908933
transform 1 0 27840 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_735
timestamp 1626908933
transform 1 0 27840 0 -1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_314
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_26
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_24
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_294
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_24
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_294
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_24
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_294
timestamp 1626908933
transform 1 0 28600 0 1 7326
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_145
timestamp 1626908933
transform 1 0 28608 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_714
timestamp 1626908933
transform 1 0 28608 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_855
timestamp 1626908933
transform 1 0 28992 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_225
timestamp 1626908933
transform 1 0 28992 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_711
timestamp 1626908933
transform 1 0 29088 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_141
timestamp 1626908933
transform 1 0 29088 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_854
timestamp 1626908933
transform 1 0 29856 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_224
timestamp 1626908933
transform 1 0 29856 0 -1 7992
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_457
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_169
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_690
timestamp 1626908933
transform 1 0 29952 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_121
timestamp 1626908933
transform 1 0 29952 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_687
timestamp 1626908933
transform 1 0 30336 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_117
timestamp 1626908933
transform 1 0 30336 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_509
timestamp 1626908933
transform 1 0 31104 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_141
timestamp 1626908933
transform 1 0 31104 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_670
timestamp 1626908933
transform 1 0 31296 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_101
timestamp 1626908933
transform 1 0 31296 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_662
timestamp 1626908933
transform 1 0 31680 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_92
timestamp 1626908933
transform 1 0 31680 0 -1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_298
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_10
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_279
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_9
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_279
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_9
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_279
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_9
timestamp 1626908933
transform 1 0 32600 0 1 7326
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_421
timestamp 1626908933
transform 1 0 32448 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_162
timestamp 1626908933
transform 1 0 32448 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_69
timestamp 1626908933
transform 1 0 32544 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_638
timestamp 1626908933
transform 1 0 32544 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_633
timestamp 1626908933
transform 1 0 32928 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_63
timestamp 1626908933
transform 1 0 32928 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_853
timestamp 1626908933
transform 1 0 33696 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_223
timestamp 1626908933
transform 1 0 33696 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_605
timestamp 1626908933
transform 1 0 33792 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_36
timestamp 1626908933
transform 1 0 33792 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_603
timestamp 1626908933
transform 1 0 34176 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_33
timestamp 1626908933
transform 1 0 34176 0 -1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_153
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_441
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_9
timestamp 1626908933
transform 1 0 34944 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_579
timestamp 1626908933
transform 1 0 34944 0 -1 7992
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1192
timestamp 1626908933
transform 1 0 144 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_404
timestamp 1626908933
transform 1 0 144 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1434
timestamp 1626908933
transform 1 0 48 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_666
timestamp 1626908933
transform 1 0 48 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1435
timestamp 1626908933
transform 1 0 240 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_667
timestamp 1626908933
transform 1 0 240 0 1 8251
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_644
timestamp 1626908933
transform 1 0 288 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_276
timestamp 1626908933
transform 1 0 288 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_420
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_161
timestamp 1626908933
transform 1 0 288 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1487
timestamp 1626908933
transform 1 0 528 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1256
timestamp 1626908933
transform 1 0 624 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_699
timestamp 1626908933
transform 1 0 528 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_468
timestamp 1626908933
transform 1 0 624 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1166
timestamp 1626908933
transform 1 0 432 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_398
timestamp 1626908933
transform 1 0 432 0 1 8325
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_137
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_425
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_398
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_128
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_398
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_128
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_398
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_128
timestamp 1626908933
transform 1 0 600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1122
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_492
timestamp 1626908933
transform 1 0 384 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1154
timestamp 1626908933
transform 1 0 816 0 1 8547
box -29 -23 29 23
use L1M1_PR  L1M1_PR_366
timestamp 1626908933
transform 1 0 816 0 1 8547
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1095
timestamp 1626908933
transform 1 0 816 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_327
timestamp 1626908933
transform 1 0 816 0 1 8103
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1186
timestamp 1626908933
transform 1 0 912 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_398
timestamp 1626908933
transform 1 0 912 0 1 8103
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_852
timestamp 1626908933
transform 1 0 1056 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_222
timestamp 1626908933
transform 1 0 1056 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_508
timestamp 1626908933
transform 1 0 864 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_140
timestamp 1626908933
transform 1 0 864 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_560
timestamp 1626908933
transform 1 0 1152 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1130
timestamp 1626908933
transform 1 0 1152 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_0
timestamp 1626908933
transform 1 0 480 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_25
timestamp 1626908933
transform 1 0 480 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_2
timestamp 1626908933
transform 1 0 864 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_11
timestamp 1626908933
transform 1 0 864 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_14
timestamp 1626908933
transform 1 0 480 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_39
timestamp 1626908933
transform 1 0 480 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_499
timestamp 1626908933
transform 1 0 1248 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_131
timestamp 1626908933
transform 1 0 1248 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1116
timestamp 1626908933
transform 1 0 1392 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_348
timestamp 1626908933
transform 1 0 1392 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_356
timestamp 1626908933
transform 1 0 1776 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1124
timestamp 1626908933
transform 1 0 1776 0 1 8399
box -32 -32 32 32
use L1M1_PR  L1M1_PR_698
timestamp 1626908933
transform 1 0 1872 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1486
timestamp 1626908933
transform 1 0 1872 0 1 8177
box -29 -23 29 23
use L1M1_PR  L1M1_PR_364
timestamp 1626908933
transform 1 0 2160 0 1 8103
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1152
timestamp 1626908933
transform 1 0 2160 0 1 8103
box -29 -23 29 23
use M1M2_PR  M1M2_PR_296
timestamp 1626908933
transform 1 0 2256 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1064
timestamp 1626908933
transform 1 0 2256 0 1 8103
box -32 -32 32 32
use M1M2_PR  M1M2_PR_347
timestamp 1626908933
transform 1 0 2256 0 1 8251
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1115
timestamp 1626908933
transform 1 0 2256 0 1 8251
box -32 -32 32 32
use L1M1_PR  L1M1_PR_456
timestamp 1626908933
transform 1 0 2064 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1244
timestamp 1626908933
transform 1 0 2064 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1066
timestamp 1626908933
transform 1 0 2064 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_298
timestamp 1626908933
transform 1 0 2064 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_498
timestamp 1626908933
transform 1 0 2208 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_130
timestamp 1626908933
transform 1 0 2208 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_23
timestamp 1626908933
transform 1 0 1920 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_48
timestamp 1626908933
transform 1 0 1920 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_559
timestamp 1626908933
transform 1 0 1440 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1129
timestamp 1626908933
transform 1 0 1440 0 -1 9324
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_264
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_534
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_264
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_534
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_264
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_534
timestamp 1626908933
transform 1 0 2600 0 1 7992
box -200 -49 200 49
use L1M1_PR  L1M1_PR_425
timestamp 1626908933
transform 1 0 2640 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1213
timestamp 1626908933
transform 1 0 2640 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_451
timestamp 1626908933
transform 1 0 2448 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1239
timestamp 1626908933
transform 1 0 2448 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_697
timestamp 1626908933
transform 1 0 2352 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1485
timestamp 1626908933
transform 1 0 2352 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_421
timestamp 1626908933
transform 1 0 2256 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1209
timestamp 1626908933
transform 1 0 2256 0 1 8251
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1167
timestamp 1626908933
transform 1 0 2640 0 1 8399
box -29 -23 29 23
use L1M1_PR  L1M1_PR_379
timestamp 1626908933
transform 1 0 2640 0 1 8399
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1129
timestamp 1626908933
transform 1 0 2400 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_499
timestamp 1626908933
transform 1 0 2400 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_412
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_153
timestamp 1626908933
transform 1 0 2496 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_273
timestamp 1626908933
transform 1 0 2688 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_641
timestamp 1626908933
transform 1 0 2688 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_493
timestamp 1626908933
transform 1 0 2880 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1123
timestamp 1626908933
transform 1 0 2880 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_351
timestamp 1626908933
transform 1 0 2832 0 1 8547
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1119
timestamp 1626908933
transform 1 0 2832 0 1 8547
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_24
timestamp 1626908933
transform 1 0 2304 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_49
timestamp 1626908933
transform 1 0 2304 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_104
timestamp 1626908933
transform 1 0 2976 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_49
timestamp 1626908933
transform 1 0 2976 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_543
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1112
timestamp 1626908933
transform 1 0 2592 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_108
timestamp 1626908933
transform 1 0 2976 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_53
timestamp 1626908933
transform 1 0 2976 0 -1 9324
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1071
timestamp 1626908933
transform 1 0 3504 0 1 8177
box -32 -32 32 32
use M1M2_PR  M1M2_PR_303
timestamp 1626908933
transform 1 0 3504 0 1 8177
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1160
timestamp 1626908933
transform 1 0 3216 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_372
timestamp 1626908933
transform 1 0 3216 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_940
timestamp 1626908933
transform 1 0 3312 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_152
timestamp 1626908933
transform 1 0 3312 0 1 8325
box -29 -23 29 23
use M1M2_PR  M1M2_PR_893
timestamp 1626908933
transform 1 0 3312 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_125
timestamp 1626908933
transform 1 0 3312 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1075
timestamp 1626908933
transform 1 0 3504 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_307
timestamp 1626908933
transform 1 0 3504 0 1 8399
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_221
timestamp 1626908933
transform 1 0 3936 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_851
timestamp 1626908933
transform 1 0 3936 0 1 7992
box -38 -49 134 715
use L1M1_PR  L1M1_PR_146
timestamp 1626908933
transform 1 0 3792 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_934
timestamp 1626908933
transform 1 0 3792 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_377
timestamp 1626908933
transform 1 0 3600 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1165
timestamp 1626908933
transform 1 0 3600 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_109
timestamp 1626908933
transform 1 0 3456 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_54
timestamp 1626908933
transform 1 0 3456 0 1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_521
timestamp 1626908933
transform 1 0 3936 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1090
timestamp 1626908933
transform 1 0 3936 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_107
timestamp 1626908933
transform 1 0 3456 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_52
timestamp 1626908933
transform 1 0 3456 0 -1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1104
timestamp 1626908933
transform 1 0 4032 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_534
timestamp 1626908933
transform 1 0 4032 0 1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_121
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_409
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_113
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_383
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_113
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_383
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_113
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_383
timestamp 1626908933
transform 1 0 4600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_160
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_419
timestamp 1626908933
transform 1 0 4992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_220
timestamp 1626908933
transform 1 0 4800 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_494
timestamp 1626908933
transform 1 0 4896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_850
timestamp 1626908933
transform 1 0 4800 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1124
timestamp 1626908933
transform 1 0 4896 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_139
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_507
timestamp 1626908933
transform 1 0 5088 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_68
timestamp 1626908933
transform 1 0 4320 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_148
timestamp 1626908933
transform 1 0 4320 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_514
timestamp 1626908933
transform 1 0 5376 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1083
timestamp 1626908933
transform 1 0 5376 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_219
timestamp 1626908933
transform 1 0 5280 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_849
timestamp 1626908933
transform 1 0 5280 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_277
timestamp 1626908933
transform 1 0 5184 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_645
timestamp 1626908933
transform 1 0 5184 0 -1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_733
timestamp 1626908933
transform 1 0 6000 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1501
timestamp 1626908933
transform 1 0 6000 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_761
timestamp 1626908933
transform 1 0 6000 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1549
timestamp 1626908933
transform 1 0 6000 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_73
timestamp 1626908933
transform 1 0 5760 0 1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_153
timestamp 1626908933
transform 1 0 5760 0 1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_78
timestamp 1626908933
transform -1 0 6240 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_158
timestamp 1626908933
transform -1 0 6240 0 -1 9324
box -38 -49 902 715
use osc_core_VIA5  osc_core_VIA5_249
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_519
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_249
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_519
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_249
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_519
timestamp 1626908933
transform 1 0 6600 0 1 7992
box -200 -49 200 49
use M1M2_PR  M1M2_PR_117
timestamp 1626908933
transform 1 0 6480 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_885
timestamp 1626908933
transform 1 0 6480 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_138
timestamp 1626908933
transform 1 0 6480 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_926
timestamp 1626908933
transform 1 0 6480 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1130
timestamp 1626908933
transform 1 0 6432 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_500
timestamp 1626908933
transform 1 0 6432 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_646
timestamp 1626908933
transform 1 0 6240 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_278
timestamp 1626908933
transform 1 0 6240 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_506
timestamp 1626908933
transform 1 0 6624 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1076
timestamp 1626908933
transform 1 0 6624 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_77
timestamp 1626908933
transform 1 0 6528 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_157
timestamp 1626908933
transform 1 0 6528 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_495
timestamp 1626908933
transform 1 0 7392 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1125
timestamp 1626908933
transform 1 0 7392 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_501
timestamp 1626908933
transform 1 0 7392 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1131
timestamp 1626908933
transform 1 0 7392 0 -1 9324
box -38 -49 134 715
use M1M2_PR  M1M2_PR_688
timestamp 1626908933
transform 1 0 7632 0 1 8325
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1456
timestamp 1626908933
transform 1 0 7632 0 1 8325
box -32 -32 32 32
use L1M1_PR  L1M1_PR_721
timestamp 1626908933
transform 1 0 7632 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1509
timestamp 1626908933
transform 1 0 7632 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_152
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_411
timestamp 1626908933
transform 1 0 7488 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_64
timestamp 1626908933
transform 1 0 7488 0 1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_144
timestamp 1626908933
transform 1 0 7488 0 1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_74
timestamp 1626908933
transform -1 0 8448 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_154
timestamp 1626908933
transform -1 0 8448 0 -1 9324
box -38 -49 902 715
use L1M1_PR  L1M1_PR_135
timestamp 1626908933
transform 1 0 8016 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_923
timestamp 1626908933
transform 1 0 8016 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_482
timestamp 1626908933
transform 1 0 8352 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1051
timestamp 1626908933
transform 1 0 8352 0 1 7992
box -38 -49 422 715
use M1M2_PR  M1M2_PR_729
timestamp 1626908933
transform 1 0 8304 0 1 8399
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1497
timestamp 1626908933
transform 1 0 8304 0 1 8399
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_393
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_105
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_368
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_98
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_368
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_98
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_368
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_98
timestamp 1626908933
transform 1 0 8600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_647
timestamp 1626908933
transform 1 0 8448 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_279
timestamp 1626908933
transform 1 0 8448 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_75
timestamp 1626908933
transform 1 0 8736 0 1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_155
timestamp 1626908933
transform 1 0 8736 0 1 7992
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_72
timestamp 1626908933
transform 1 0 8640 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_152
timestamp 1626908933
transform 1 0 8640 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1035
timestamp 1626908933
transform 1 0 9504 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_466
timestamp 1626908933
transform 1 0 9504 0 -1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1540
timestamp 1626908933
transform 1 0 8880 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_911
timestamp 1626908933
transform 1 0 9264 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_752
timestamp 1626908933
transform 1 0 8880 0 1 8325
box -29 -23 29 23
use L1M1_PR  L1M1_PR_123
timestamp 1626908933
transform 1 0 9264 0 1 8325
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1023
timestamp 1626908933
transform 1 0 9600 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_454
timestamp 1626908933
transform 1 0 9600 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_159
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_418
timestamp 1626908933
transform 1 0 9984 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_447
timestamp 1626908933
transform 1 0 10080 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1016
timestamp 1626908933
transform 1 0 10080 0 1 7992
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_234
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_504
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_234
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_504
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_234
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_504
timestamp 1626908933
transform 1 0 10600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_462
timestamp 1626908933
transform 1 0 10464 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1032
timestamp 1626908933
transform 1 0 10464 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_67
timestamp 1626908933
transform -1 0 10752 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_147
timestamp 1626908933
transform -1 0 10752 0 -1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_129
timestamp 1626908933
transform 1 0 10752 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_497
timestamp 1626908933
transform 1 0 10752 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_205
timestamp 1626908933
transform 1 0 10944 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_835
timestamp 1626908933
transform 1 0 10944 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_424
timestamp 1626908933
transform 1 0 11328 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_993
timestamp 1626908933
transform 1 0 11328 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_218
timestamp 1626908933
transform 1 0 11232 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_848
timestamp 1626908933
transform 1 0 11232 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_455
timestamp 1626908933
transform 1 0 11040 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1025
timestamp 1626908933
transform 1 0 11040 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_204
timestamp 1626908933
transform 1 0 12000 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_834
timestamp 1626908933
transform 1 0 12000 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_128
timestamp 1626908933
transform 1 0 11808 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_496
timestamp 1626908933
transform 1 0 11808 0 -1 9324
box -38 -49 230 715
use osc_core_VIA4  osc_core_VIA4_377
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_89
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_353
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_83
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_353
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_83
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_353
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_83
timestamp 1626908933
transform 1 0 12600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_988
timestamp 1626908933
transform 1 0 12096 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_419
timestamp 1626908933
transform 1 0 12096 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_441
timestamp 1626908933
transform 1 0 11712 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1011
timestamp 1626908933
transform 1 0 11712 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_217
timestamp 1626908933
transform 1 0 12864 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_847
timestamp 1626908933
transform 1 0 12864 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_151
timestamp 1626908933
transform 1 0 12480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_410
timestamp 1626908933
transform 1 0 12480 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_427
timestamp 1626908933
transform 1 0 12960 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_997
timestamp 1626908933
transform 1 0 12960 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_406
timestamp 1626908933
transform 1 0 12480 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_975
timestamp 1626908933
transform 1 0 12480 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_426
timestamp 1626908933
transform 1 0 12960 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_996
timestamp 1626908933
transform 1 0 12960 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_397
timestamp 1626908933
transform 1 0 12576 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_966
timestamp 1626908933
transform 1 0 12576 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_943
timestamp 1626908933
transform 1 0 13920 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_374
timestamp 1626908933
transform 1 0 13920 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_495
timestamp 1626908933
transform 1 0 13728 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_127
timestamp 1626908933
transform 1 0 13728 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_846
timestamp 1626908933
transform 1 0 13728 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_216
timestamp 1626908933
transform 1 0 13728 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_944
timestamp 1626908933
transform 1 0 13824 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_375
timestamp 1626908933
transform 1 0 13824 0 1 7992
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_219
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_489
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_219
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_489
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_219
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_489
timestamp 1626908933
transform 1 0 14600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_158
timestamp 1626908933
transform 1 0 14976 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_417
timestamp 1626908933
transform 1 0 14976 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_413
timestamp 1626908933
transform 1 0 14208 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_983
timestamp 1626908933
transform 1 0 14208 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_412
timestamp 1626908933
transform 1 0 14304 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_982
timestamp 1626908933
transform 1 0 14304 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_833
timestamp 1626908933
transform 1 0 15072 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_203
timestamp 1626908933
transform 1 0 15072 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_924
timestamp 1626908933
transform 1 0 15168 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_355
timestamp 1626908933
transform 1 0 15168 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_845
timestamp 1626908933
transform 1 0 15072 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_215
timestamp 1626908933
transform 1 0 15072 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_925
timestamp 1626908933
transform 1 0 15168 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_356
timestamp 1626908933
transform 1 0 15168 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_962
timestamp 1626908933
transform 1 0 15552 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_392
timestamp 1626908933
transform 1 0 15552 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_963
timestamp 1626908933
transform 1 0 15552 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_393
timestamp 1626908933
transform 1 0 15552 0 1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_361
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_73
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_338
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_68
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_338
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_68
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_338
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_68
timestamp 1626908933
transform 1 0 16600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_506
timestamp 1626908933
transform 1 0 16320 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_138
timestamp 1626908933
transform 1 0 16320 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_331
timestamp 1626908933
transform 1 0 16512 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_900
timestamp 1626908933
transform 1 0 16512 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_367
timestamp 1626908933
transform 1 0 16896 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_937
timestamp 1626908933
transform 1 0 16896 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_330
timestamp 1626908933
transform 1 0 16320 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_899
timestamp 1626908933
transform 1 0 16320 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_366
timestamp 1626908933
transform 1 0 16704 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_936
timestamp 1626908933
transform 1 0 16704 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_214
timestamp 1626908933
transform 1 0 17664 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_844
timestamp 1626908933
transform 1 0 17664 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_126
timestamp 1626908933
transform 1 0 17568 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_494
timestamp 1626908933
transform 1 0 17568 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_150
timestamp 1626908933
transform 1 0 17472 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_409
timestamp 1626908933
transform 1 0 17472 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_306
timestamp 1626908933
transform 1 0 17760 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_875
timestamp 1626908933
transform 1 0 17760 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_305
timestamp 1626908933
transform 1 0 17760 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_874
timestamp 1626908933
transform 1 0 17760 0 -1 9324
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_204
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_474
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_204
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_474
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_204
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_474
timestamp 1626908933
transform 1 0 18600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_344
timestamp 1626908933
transform 1 0 18144 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_914
timestamp 1626908933
transform 1 0 18144 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_343
timestamp 1626908933
transform 1 0 18144 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_913
timestamp 1626908933
transform 1 0 18144 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_137
timestamp 1626908933
transform 1 0 18912 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_505
timestamp 1626908933
transform 1 0 18912 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_213
timestamp 1626908933
transform 1 0 19104 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_843
timestamp 1626908933
transform 1 0 19104 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_202
timestamp 1626908933
transform 1 0 19296 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_832
timestamp 1626908933
transform 1 0 19296 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_322
timestamp 1626908933
transform 1 0 19200 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_892
timestamp 1626908933
transform 1 0 19200 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_321
timestamp 1626908933
transform 1 0 19392 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_891
timestamp 1626908933
transform 1 0 19392 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_286
timestamp 1626908933
transform 1 0 18912 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_855
timestamp 1626908933
transform 1 0 18912 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_157
timestamp 1626908933
transform 1 0 19968 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_416
timestamp 1626908933
transform 1 0 19968 0 1 7992
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_323
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_53
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_323
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_53
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_323
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_53
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_57
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_345
timestamp 1626908933
transform 1 0 20600 0 1 8658
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_493
timestamp 1626908933
transform 1 0 20160 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_125
timestamp 1626908933
transform 1 0 20160 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_303
timestamp 1626908933
transform 1 0 20064 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_873
timestamp 1626908933
transform 1 0 20064 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_270
timestamp 1626908933
transform 1 0 20352 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_839
timestamp 1626908933
transform 1 0 20352 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_861
timestamp 1626908933
transform 1 0 20736 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_291
timestamp 1626908933
transform 1 0 20736 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_492
timestamp 1626908933
transform 1 0 21504 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_124
timestamp 1626908933
transform 1 0 21504 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_504
timestamp 1626908933
transform 1 0 20832 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_136
timestamp 1626908933
transform 1 0 20832 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_824
timestamp 1626908933
transform 1 0 21024 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_255
timestamp 1626908933
transform 1 0 21024 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_847
timestamp 1626908933
transform 1 0 21408 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_277
timestamp 1626908933
transform 1 0 21408 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_212
timestamp 1626908933
transform 1 0 22176 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_842
timestamp 1626908933
transform 1 0 22176 0 1 7992
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_189
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_459
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_189
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_459
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_189
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_459
timestamp 1626908933
transform 1 0 22600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_236
timestamp 1626908933
transform 1 0 22272 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_805
timestamp 1626908933
transform 1 0 22272 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_267
timestamp 1626908933
transform 1 0 21696 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_837
timestamp 1626908933
transform 1 0 21696 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_831
timestamp 1626908933
transform 1 0 22560 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_201
timestamp 1626908933
transform 1 0 22560 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_821
timestamp 1626908933
transform 1 0 22656 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_251
timestamp 1626908933
transform 1 0 22656 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_408
timestamp 1626908933
transform 1 0 22464 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_149
timestamp 1626908933
transform 1 0 22464 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_822
timestamp 1626908933
transform 1 0 22656 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_252
timestamp 1626908933
transform 1 0 22656 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_786
timestamp 1626908933
transform 1 0 23424 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_217
timestamp 1626908933
transform 1 0 23424 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_787
timestamp 1626908933
transform 1 0 23424 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_218
timestamp 1626908933
transform 1 0 23424 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_830
timestamp 1626908933
transform 1 0 23808 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_200
timestamp 1626908933
transform 1 0 23808 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_798
timestamp 1626908933
transform 1 0 23904 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_228
timestamp 1626908933
transform 1 0 23904 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_841
timestamp 1626908933
transform 1 0 23808 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_211
timestamp 1626908933
transform 1 0 23808 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_799
timestamp 1626908933
transform 1 0 23904 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_229
timestamp 1626908933
transform 1 0 23904 0 1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_329
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_41
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_308
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_38
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_308
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_38
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_308
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_38
timestamp 1626908933
transform 1 0 24600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_491
timestamp 1626908933
transform 1 0 24672 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_123
timestamp 1626908933
transform 1 0 24672 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_642
timestamp 1626908933
transform 1 0 24672 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_274
timestamp 1626908933
transform 1 0 24672 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_496
timestamp 1626908933
transform 1 0 24864 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1126
timestamp 1626908933
transform 1 0 24864 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_156
timestamp 1626908933
transform 1 0 24960 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_415
timestamp 1626908933
transform 1 0 24960 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_135
timestamp 1626908933
transform 1 0 25056 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_503
timestamp 1626908933
transform 1 0 25056 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_200
timestamp 1626908933
transform 1 0 24864 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_769
timestamp 1626908933
transform 1 0 24864 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_777
timestamp 1626908933
transform 1 0 25248 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_207
timestamp 1626908933
transform 1 0 25248 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_749
timestamp 1626908933
transform 1 0 26016 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_180
timestamp 1626908933
transform 1 0 26016 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_778
timestamp 1626908933
transform 1 0 25248 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_208
timestamp 1626908933
transform 1 0 25248 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_750
timestamp 1626908933
transform 1 0 26016 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_181
timestamp 1626908933
transform 1 0 26016 0 1 7992
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_444
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_174
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_444
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_174
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_444
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_174
timestamp 1626908933
transform 1 0 26600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_829
timestamp 1626908933
transform 1 0 26400 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_199
timestamp 1626908933
transform 1 0 26400 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_840
timestamp 1626908933
transform 1 0 26400 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_210
timestamp 1626908933
transform 1 0 26400 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_186
timestamp 1626908933
transform 1 0 26496 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_756
timestamp 1626908933
transform 1 0 26496 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_185
timestamp 1626908933
transform 1 0 26496 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_755
timestamp 1626908933
transform 1 0 26496 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_828
timestamp 1626908933
transform 1 0 27264 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_198
timestamp 1626908933
transform 1 0 27264 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1132
timestamp 1626908933
transform 1 0 27360 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_502
timestamp 1626908933
transform 1 0 27360 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_407
timestamp 1626908933
transform 1 0 27456 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_148
timestamp 1626908933
transform 1 0 27456 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_490
timestamp 1626908933
transform 1 0 27552 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_122
timestamp 1626908933
transform 1 0 27552 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_502
timestamp 1626908933
transform 1 0 27264 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_134
timestamp 1626908933
transform 1 0 27264 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_197
timestamp 1626908933
transform 1 0 27744 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_827
timestamp 1626908933
transform 1 0 27744 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_163
timestamp 1626908933
transform 1 0 27456 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_732
timestamp 1626908933
transform 1 0 27456 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_164
timestamp 1626908933
transform 1 0 27840 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_734
timestamp 1626908933
transform 1 0 27840 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_163
timestamp 1626908933
transform 1 0 27840 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_733
timestamp 1626908933
transform 1 0 27840 0 -1 9324
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_313
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_25
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_23
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_293
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_23
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_293
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_23
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_293
timestamp 1626908933
transform 1 0 28600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_144
timestamp 1626908933
transform 1 0 28608 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_713
timestamp 1626908933
transform 1 0 28608 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_143
timestamp 1626908933
transform 1 0 28608 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_712
timestamp 1626908933
transform 1 0 28608 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_826
timestamp 1626908933
transform 1 0 28992 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_196
timestamp 1626908933
transform 1 0 28992 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_839
timestamp 1626908933
transform 1 0 28992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_209
timestamp 1626908933
transform 1 0 28992 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_709
timestamp 1626908933
transform 1 0 29088 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_139
timestamp 1626908933
transform 1 0 29088 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_825
timestamp 1626908933
transform 1 0 29856 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_195
timestamp 1626908933
transform 1 0 29856 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_710
timestamp 1626908933
transform 1 0 29088 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_140
timestamp 1626908933
transform 1 0 29088 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1127
timestamp 1626908933
transform 1 0 29856 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_497
timestamp 1626908933
transform 1 0 29856 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_208
timestamp 1626908933
transform 1 0 30240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_838
timestamp 1626908933
transform 1 0 30240 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_155
timestamp 1626908933
transform 1 0 29952 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_414
timestamp 1626908933
transform 1 0 29952 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_133
timestamp 1626908933
transform 1 0 30048 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_501
timestamp 1626908933
transform 1 0 30048 0 1 7992
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_159
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_429
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_159
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_429
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_159
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_429
timestamp 1626908933
transform 1 0 30600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_116
timestamp 1626908933
transform 1 0 30336 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_686
timestamp 1626908933
transform 1 0 30336 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_115
timestamp 1626908933
transform 1 0 30336 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_685
timestamp 1626908933
transform 1 0 30336 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_120
timestamp 1626908933
transform 1 0 29952 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_689
timestamp 1626908933
transform 1 0 29952 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_489
timestamp 1626908933
transform 1 0 31104 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_121
timestamp 1626908933
transform 1 0 31104 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_668
timestamp 1626908933
transform 1 0 31296 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_99
timestamp 1626908933
transform 1 0 31296 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_500
timestamp 1626908933
transform 1 0 31104 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_132
timestamp 1626908933
transform 1 0 31104 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_669
timestamp 1626908933
transform 1 0 31296 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_100
timestamp 1626908933
transform 1 0 31296 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_660
timestamp 1626908933
transform 1 0 31680 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_90
timestamp 1626908933
transform 1 0 31680 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_661
timestamp 1626908933
transform 1 0 31680 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_91
timestamp 1626908933
transform 1 0 31680 0 1 7992
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_297
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_9
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_278
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_8
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_278
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_8
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_278
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_8
timestamp 1626908933
transform 1 0 32600 0 1 8658
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_406
timestamp 1626908933
transform 1 0 32448 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_147
timestamp 1626908933
transform 1 0 32448 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_837
timestamp 1626908933
transform 1 0 32448 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_207
timestamp 1626908933
transform 1 0 32448 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_68
timestamp 1626908933
transform 1 0 32544 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_637
timestamp 1626908933
transform 1 0 32544 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_67
timestamp 1626908933
transform 1 0 32544 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_636
timestamp 1626908933
transform 1 0 32544 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_631
timestamp 1626908933
transform 1 0 32928 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_61
timestamp 1626908933
transform 1 0 32928 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_632
timestamp 1626908933
transform 1 0 32928 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_62
timestamp 1626908933
transform 1 0 32928 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_206
timestamp 1626908933
transform 1 0 33696 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_836
timestamp 1626908933
transform 1 0 33696 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_194
timestamp 1626908933
transform 1 0 33696 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_824
timestamp 1626908933
transform 1 0 33696 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_32
timestamp 1626908933
transform 1 0 34176 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_602
timestamp 1626908933
transform 1 0 34176 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_35
timestamp 1626908933
transform 1 0 33792 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_604
timestamp 1626908933
transform 1 0 33792 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_31
timestamp 1626908933
transform 1 0 34176 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_601
timestamp 1626908933
transform 1 0 34176 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_34
timestamp 1626908933
transform 1 0 33792 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_603
timestamp 1626908933
transform 1 0 33792 0 -1 9324
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_414
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_144
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_414
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_144
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_414
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_144
timestamp 1626908933
transform 1 0 34600 0 1 7992
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_578
timestamp 1626908933
transform 1 0 34944 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_8
timestamp 1626908933
transform 1 0 34944 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_643
timestamp 1626908933
transform 1 0 35424 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_275
timestamp 1626908933
transform 1 0 35424 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_578
timestamp 1626908933
transform 1 0 35040 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_9
timestamp 1626908933
transform 1 0 35040 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_413
timestamp 1626908933
transform 1 0 34944 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_154
timestamp 1626908933
transform 1 0 34944 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1128
timestamp 1626908933
transform 1 0 35616 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_498
timestamp 1626908933
transform 1 0 35616 0 1 7992
box -38 -49 134 715
use M1M2_PR  M1M2_PR_665
timestamp 1626908933
transform 1 0 144 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1433
timestamp 1626908933
transform 1 0 144 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_400
timestamp 1626908933
transform 1 0 336 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1168
timestamp 1626908933
transform 1 0 336 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_696
timestamp 1626908933
transform 1 0 432 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1484
timestamp 1626908933
transform 1 0 432 0 1 8769
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_146
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_405
timestamp 1626908933
transform 1 0 288 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_503
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1133
timestamp 1626908933
transform 1 0 384 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_13
timestamp 1626908933
transform 1 0 480 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_38
timestamp 1626908933
transform 1 0 480 0 1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_415
timestamp 1626908933
transform 1 0 912 0 1 8769
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1203
timestamp 1626908933
transform 1 0 912 0 1 8769
box -29 -23 29 23
use M1M2_PR  M1M2_PR_394
timestamp 1626908933
transform 1 0 624 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1162
timestamp 1626908933
transform 1 0 624 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_467
timestamp 1626908933
transform 1 0 624 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1255
timestamp 1626908933
transform 1 0 624 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_305
timestamp 1626908933
transform 1 0 720 0 1 9213
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1093
timestamp 1626908933
transform 1 0 720 0 1 9213
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_556
timestamp 1626908933
transform 1 0 864 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1125
timestamp 1626908933
transform 1 0 864 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_488
timestamp 1626908933
transform 1 0 1248 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_120
timestamp 1626908933
transform 1 0 1248 0 1 9324
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1108
timestamp 1626908933
transform 1 0 1008 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1106
timestamp 1626908933
transform 1 0 1296 0 1 8843
box -32 -32 32 32
use M1M2_PR  M1M2_PR_340
timestamp 1626908933
transform 1 0 1008 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_338
timestamp 1626908933
transform 1 0 1296 0 1 8843
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1128
timestamp 1626908933
transform 1 0 1440 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_558
timestamp 1626908933
transform 1 0 1440 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1116
timestamp 1626908933
transform 1 0 2208 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_546
timestamp 1626908933
transform 1 0 2208 0 1 9324
box -38 -49 806 715
use L1M1_PR  L1M1_PR_378
timestamp 1626908933
transform 1 0 3216 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1166
timestamp 1626908933
transform 1 0 3216 0 1 8991
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_568
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_280
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_263
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_533
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_263
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_533
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_263
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_533
timestamp 1626908933
transform 1 0 2600 0 1 9324
box -200 -49 200 49
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_55
timestamp 1626908933
transform 1 0 2976 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_0
timestamp 1626908933
transform 1 0 2976 0 1 9324
box -38 -49 518 715
use L1M1_PR  L1M1_PR_939
timestamp 1626908933
transform 1 0 3312 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_151
timestamp 1626908933
transform 1 0 3312 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_892
timestamp 1626908933
transform 1 0 3312 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_124
timestamp 1626908933
transform 1 0 3312 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1074
timestamp 1626908933
transform 1 0 3504 0 1 8917
box -32 -32 32 32
use M1M2_PR  M1M2_PR_306
timestamp 1626908933
transform 1 0 3504 0 1 8917
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1164
timestamp 1626908933
transform 1 0 3600 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_376
timestamp 1626908933
transform 1 0 3600 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1016
timestamp 1626908933
transform 1 0 3696 0 1 9213
box -32 -32 32 32
use M1M2_PR  M1M2_PR_248
timestamp 1626908933
transform 1 0 3696 0 1 9213
box -32 -32 32 32
use L1M1_PR  L1M1_PR_145
timestamp 1626908933
transform 1 0 3792 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_933
timestamp 1626908933
transform 1 0 3792 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_280
timestamp 1626908933
transform 1 0 3936 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_648
timestamp 1626908933
transform 1 0 3936 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_12
timestamp 1626908933
transform -1 0 4992 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_92
timestamp 1626908933
transform -1 0 4992 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_106
timestamp 1626908933
transform 1 0 3456 0 1 9324
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_51
timestamp 1626908933
transform 1 0 3456 0 1 9324
box -38 -49 518 715
use M1M2_PR  M1M2_PR_709
timestamp 1626908933
transform 1 0 4272 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1477
timestamp 1626908933
transform 1 0 4272 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_738
timestamp 1626908933
transform 1 0 4464 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1526
timestamp 1626908933
transform 1 0 4464 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_710
timestamp 1626908933
transform 1 0 4272 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1478
timestamp 1626908933
transform 1 0 4272 0 1 8769
box -32 -32 32 32
use L1M1_PR  L1M1_PR_143
timestamp 1626908933
transform 1 0 4848 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_931
timestamp 1626908933
transform 1 0 4848 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_145
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_404
timestamp 1626908933
transform 1 0 4992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_521
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1091
timestamp 1626908933
transform 1 0 5088 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_94
timestamp 1626908933
transform 1 0 5856 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_14
timestamp 1626908933
transform 1 0 5856 0 1 9324
box -38 -49 902 715
use M1M2_PR  M1M2_PR_1513
timestamp 1626908933
transform 1 0 6000 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_745
timestamp 1626908933
transform 1 0 6000 0 1 8991
box -32 -32 32 32
use L1M1_PR  L1M1_PR_930
timestamp 1626908933
transform 1 0 5520 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_142
timestamp 1626908933
transform 1 0 5520 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1557
timestamp 1626908933
transform 1 0 6096 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_769
timestamp 1626908933
transform 1 0 6096 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_116
timestamp 1626908933
transform 1 0 6480 0 1 9065
box -32 -32 32 32
use M1M2_PR  M1M2_PR_884
timestamp 1626908933
transform 1 0 6480 0 1 9065
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_248
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_518
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_248
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_518
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_248
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_518
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_552
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_264
timestamp 1626908933
transform 1 0 6600 0 1 9324
box -200 -142 200 178
use L1M1_PR  L1M1_PR_764
timestamp 1626908933
transform 1 0 6672 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1552
timestamp 1626908933
transform 1 0 6672 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_494
timestamp 1626908933
transform 1 0 6912 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1063
timestamp 1626908933
transform 1 0 6912 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_119
timestamp 1626908933
transform 1 0 6720 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_487
timestamp 1626908933
transform 1 0 6720 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_145
timestamp 1626908933
transform 1 0 7392 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_65
timestamp 1626908933
transform 1 0 7392 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1134
timestamp 1626908933
transform 1 0 7296 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_504
timestamp 1626908933
transform 1 0 7296 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_925
timestamp 1626908933
transform 1 0 7056 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_137
timestamp 1626908933
transform 1 0 7056 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_924
timestamp 1626908933
transform 1 0 7728 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_136
timestamp 1626908933
transform 1 0 7728 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1545
timestamp 1626908933
transform 1 0 8304 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_757
timestamp 1626908933
transform 1 0 8304 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1496
timestamp 1626908933
transform 1 0 8304 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_728
timestamp 1626908933
transform 1 0 8304 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1474
timestamp 1626908933
transform 1 0 7920 0 1 8769
box -32 -32 32 32
use M1M2_PR  M1M2_PR_706
timestamp 1626908933
transform 1 0 7920 0 1 8769
box -32 -32 32 32
use M3M4_PR  M3M4_PR_32
timestamp 1626908933
transform 1 0 8112 0 1 9431
box -38 -33 38 33
use M3M4_PR  M3M4_PR_11
timestamp 1626908933
transform 1 0 8112 0 1 9431
box -38 -33 38 33
use M2M3_PR  M2M3_PR_71
timestamp 1626908933
transform 1 0 8112 0 1 9431
box -33 -37 33 37
use M2M3_PR  M2M3_PR_12
timestamp 1626908933
transform 1 0 8112 0 1 9431
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_649
timestamp 1626908933
transform 1 0 8256 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_281
timestamp 1626908933
transform 1 0 8256 0 1 9324
box -38 -49 230 715
use L1M1_PR  L1M1_PR_753
timestamp 1626908933
transform 1 0 8784 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1541
timestamp 1626908933
transform 1 0 8784 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_505
timestamp 1626908933
transform 1 0 8448 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1135
timestamp 1626908933
transform 1 0 8448 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_71
timestamp 1626908933
transform 1 0 8544 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_151
timestamp 1626908933
transform 1 0 8544 0 1 9324
box -38 -49 902 715
use M2M3_PR  M2M3_PR_65
timestamp 1626908933
transform 1 0 9072 0 1 9431
box -33 -37 33 37
use M2M3_PR  M2M3_PR_6
timestamp 1626908933
transform 1 0 9072 0 1 9431
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_823
timestamp 1626908933
transform 1 0 9408 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_193
timestamp 1626908933
transform 1 0 9408 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1034
timestamp 1626908933
transform 1 0 9504 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_465
timestamp 1626908933
transform 1 0 9504 0 1 9324
box -38 -49 422 715
use L1M1_PR  L1M1_PR_910
timestamp 1626908933
transform 1 0 9360 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_122
timestamp 1626908933
transform 1 0 9360 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_121
timestamp 1626908933
transform 1 0 10032 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_909
timestamp 1626908933
transform 1 0 10032 0 1 8991
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_144
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_403
timestamp 1626908933
transform 1 0 9984 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_191
timestamp 1626908933
transform 1 0 10080 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_192
timestamp 1626908933
transform 1 0 9888 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_821
timestamp 1626908933
transform 1 0 10080 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_822
timestamp 1626908933
transform 1 0 9888 0 1 9324
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1505
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -29 -23 29 23
use L1M1_PR  L1M1_PR_717
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1454
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -32 -32 32 32
use M1M2_PR  M1M2_PR_686
timestamp 1626908933
transform 1 0 10320 0 1 8991
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_503
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_233
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_503
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_233
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_503
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_233
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_248
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_536
timestamp 1626908933
transform 1 0 10600 0 1 9324
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_461
timestamp 1626908933
transform 1 0 10176 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1031
timestamp 1626908933
transform 1 0 10176 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_84
timestamp 1626908933
transform 1 0 10944 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_4
timestamp 1626908933
transform 1 0 10944 0 1 9324
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_486
timestamp 1626908933
transform 1 0 11808 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_118
timestamp 1626908933
transform 1 0 11808 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_987
timestamp 1626908933
transform 1 0 12000 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_418
timestamp 1626908933
transform 1 0 12000 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1010
timestamp 1626908933
transform 1 0 12384 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_440
timestamp 1626908933
transform 1 0 12384 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_820
timestamp 1626908933
transform 1 0 13152 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_190
timestamp 1626908933
transform 1 0 13152 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_956
timestamp 1626908933
transform 1 0 13248 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_387
timestamp 1626908933
transform 1 0 13248 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_994
timestamp 1626908933
transform 1 0 13632 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_424
timestamp 1626908933
transform 1 0 13632 0 1 9324
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_520
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_232
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_218
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_488
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_218
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_488
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_218
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_488
timestamp 1626908933
transform 1 0 14600 0 1 9324
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_143
timestamp 1626908933
transform 1 0 14976 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_402
timestamp 1626908933
transform 1 0 14976 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_189
timestamp 1626908933
transform 1 0 14784 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_506
timestamp 1626908933
transform 1 0 14880 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_819
timestamp 1626908933
transform 1 0 14784 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1136
timestamp 1626908933
transform 1 0 14880 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_370
timestamp 1626908933
transform 1 0 14400 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_939
timestamp 1626908933
transform 1 0 14400 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_923
timestamp 1626908933
transform 1 0 15168 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_354
timestamp 1626908933
transform 1 0 15168 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_818
timestamp 1626908933
transform 1 0 15072 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_188
timestamp 1626908933
transform 1 0 15072 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_961
timestamp 1626908933
transform 1 0 15552 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_391
timestamp 1626908933
transform 1 0 15552 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_935
timestamp 1626908933
transform 1 0 16896 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_365
timestamp 1626908933
transform 1 0 16896 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_485
timestamp 1626908933
transform 1 0 16320 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_117
timestamp 1626908933
transform 1 0 16320 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_898
timestamp 1626908933
transform 1 0 16512 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_329
timestamp 1626908933
transform 1 0 16512 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_817
timestamp 1626908933
transform 1 0 17664 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_187
timestamp 1626908933
transform 1 0 17664 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_873
timestamp 1626908933
transform 1 0 17760 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_304
timestamp 1626908933
transform 1 0 17760 0 1 9324
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_504
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_216
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_203
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_473
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_203
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_473
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_203
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_473
timestamp 1626908933
transform 1 0 18600 0 1 9324
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_342
timestamp 1626908933
transform 1 0 18144 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_912
timestamp 1626908933
transform 1 0 18144 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_816
timestamp 1626908933
transform 1 0 19104 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_186
timestamp 1626908933
transform 1 0 19104 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_484
timestamp 1626908933
transform 1 0 18912 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_116
timestamp 1626908933
transform 1 0 18912 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_890
timestamp 1626908933
transform 1 0 19200 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_320
timestamp 1626908933
transform 1 0 19200 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_872
timestamp 1626908933
transform 1 0 20064 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_302
timestamp 1626908933
transform 1 0 20064 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_401
timestamp 1626908933
transform 1 0 19968 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_142
timestamp 1626908933
transform 1 0 19968 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_483
timestamp 1626908933
transform 1 0 20832 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_115
timestamp 1626908933
transform 1 0 20832 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_823
timestamp 1626908933
transform 1 0 21024 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_254
timestamp 1626908933
transform 1 0 21024 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_846
timestamp 1626908933
transform 1 0 21408 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_276
timestamp 1626908933
transform 1 0 21408 0 1 9324
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_488
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_200
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_458
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_188
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_458
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_188
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_458
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_188
timestamp 1626908933
transform 1 0 22600 0 1 9324
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_815
timestamp 1626908933
transform 1 0 22176 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_185
timestamp 1626908933
transform 1 0 22176 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_235
timestamp 1626908933
transform 1 0 22272 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_804
timestamp 1626908933
transform 1 0 22272 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_820
timestamp 1626908933
transform 1 0 22656 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_250
timestamp 1626908933
transform 1 0 22656 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_785
timestamp 1626908933
transform 1 0 23424 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_216
timestamp 1626908933
transform 1 0 23424 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_814
timestamp 1626908933
transform 1 0 23808 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_184
timestamp 1626908933
transform 1 0 23808 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_797
timestamp 1626908933
transform 1 0 23904 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_227
timestamp 1626908933
transform 1 0 23904 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_482
timestamp 1626908933
transform 1 0 25056 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_114
timestamp 1626908933
transform 1 0 25056 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_400
timestamp 1626908933
transform 1 0 24960 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_141
timestamp 1626908933
transform 1 0 24960 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_650
timestamp 1626908933
transform 1 0 24672 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_282
timestamp 1626908933
transform 1 0 24672 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1137
timestamp 1626908933
transform 1 0 24864 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_507
timestamp 1626908933
transform 1 0 24864 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_776
timestamp 1626908933
transform 1 0 25248 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_206
timestamp 1626908933
transform 1 0 25248 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_748
timestamp 1626908933
transform 1 0 26016 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_179
timestamp 1626908933
transform 1 0 26016 0 1 9324
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_472
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_184
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_443
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_173
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_443
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_173
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_443
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_173
timestamp 1626908933
transform 1 0 26600 0 1 9324
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_813
timestamp 1626908933
transform 1 0 26400 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_183
timestamp 1626908933
transform 1 0 26400 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_184
timestamp 1626908933
transform 1 0 26496 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_754
timestamp 1626908933
transform 1 0 26496 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_113
timestamp 1626908933
transform 1 0 27552 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_481
timestamp 1626908933
transform 1 0 27552 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_140
timestamp 1626908933
transform 1 0 27456 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_399
timestamp 1626908933
transform 1 0 27456 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_182
timestamp 1626908933
transform 1 0 27264 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_508
timestamp 1626908933
transform 1 0 27360 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_812
timestamp 1626908933
transform 1 0 27264 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1138
timestamp 1626908933
transform 1 0 27360 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_181
timestamp 1626908933
transform 1 0 27744 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_811
timestamp 1626908933
transform 1 0 27744 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_162
timestamp 1626908933
transform 1 0 27840 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_732
timestamp 1626908933
transform 1 0 27840 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_711
timestamp 1626908933
transform 1 0 28608 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_142
timestamp 1626908933
transform 1 0 28608 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_810
timestamp 1626908933
transform 1 0 28992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_180
timestamp 1626908933
transform 1 0 28992 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_708
timestamp 1626908933
transform 1 0 29088 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_138
timestamp 1626908933
transform 1 0 29088 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1139
timestamp 1626908933
transform 1 0 29856 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_509
timestamp 1626908933
transform 1 0 29856 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_179
timestamp 1626908933
transform 1 0 30240 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_809
timestamp 1626908933
transform 1 0 30240 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_139
timestamp 1626908933
transform 1 0 29952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_398
timestamp 1626908933
transform 1 0 29952 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_112
timestamp 1626908933
transform 1 0 30048 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_480
timestamp 1626908933
transform 1 0 30048 0 1 9324
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_158
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_428
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_158
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_428
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_158
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_428
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_168
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_456
timestamp 1626908933
transform 1 0 30600 0 1 9324
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_114
timestamp 1626908933
transform 1 0 30336 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_684
timestamp 1626908933
transform 1 0 30336 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_479
timestamp 1626908933
transform 1 0 31104 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_111
timestamp 1626908933
transform 1 0 31104 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_667
timestamp 1626908933
transform 1 0 31296 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_98
timestamp 1626908933
transform 1 0 31296 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_659
timestamp 1626908933
transform 1 0 31680 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_89
timestamp 1626908933
transform 1 0 31680 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_808
timestamp 1626908933
transform 1 0 32448 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_178
timestamp 1626908933
transform 1 0 32448 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_635
timestamp 1626908933
transform 1 0 32544 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_66
timestamp 1626908933
transform 1 0 32544 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_630
timestamp 1626908933
transform 1 0 32928 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_60
timestamp 1626908933
transform 1 0 32928 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_807
timestamp 1626908933
transform 1 0 33696 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_177
timestamp 1626908933
transform 1 0 33696 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_602
timestamp 1626908933
transform 1 0 33792 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_33
timestamp 1626908933
transform 1 0 33792 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_600
timestamp 1626908933
transform 1 0 34176 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_30
timestamp 1626908933
transform 1 0 34176 0 1 9324
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_413
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_143
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_413
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_143
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_413
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_143
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_152
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_440
timestamp 1626908933
transform 1 0 34600 0 1 9324
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_138
timestamp 1626908933
transform 1 0 34944 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_397
timestamp 1626908933
transform 1 0 34944 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_8
timestamp 1626908933
transform 1 0 35040 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_577
timestamp 1626908933
transform 1 0 35040 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_283
timestamp 1626908933
transform 1 0 35424 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_651
timestamp 1626908933
transform 1 0 35424 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_510
timestamp 1626908933
transform 1 0 35616 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1140
timestamp 1626908933
transform 1 0 35616 0 1 9324
box -38 -49 134 715
use M2M3_PR  M2M3_PR_107
timestamp 1626908933
transform 1 0 48 0 1 10163
box -33 -37 33 37
use M2M3_PR  M2M3_PR_48
timestamp 1626908933
transform 1 0 48 0 1 10163
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1141
timestamp 1626908933
transform 1 0 288 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_511
timestamp 1626908933
transform 1 0 288 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1432
timestamp 1626908933
transform 1 0 48 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_664
timestamp 1626908933
transform 1 0 48 0 1 9509
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1483
timestamp 1626908933
transform 1 0 528 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_695
timestamp 1626908933
transform 1 0 528 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1196
timestamp 1626908933
transform 1 0 816 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_408
timestamp 1626908933
transform 1 0 816 0 1 9583
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1254
timestamp 1626908933
transform 1 0 624 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_466
timestamp 1626908933
transform 1 0 624 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1161
timestamp 1626908933
transform 1 0 624 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_393
timestamp 1626908933
transform 1 0 624 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1088
timestamp 1626908933
transform 1 0 816 0 1 9805
box -29 -23 29 23
use L1M1_PR  L1M1_PR_300
timestamp 1626908933
transform 1 0 816 0 1 9805
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_397
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_127
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_397
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_127
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_397
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_127
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1187
timestamp 1626908933
transform 1 0 816 0 1 10175
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1085
timestamp 1626908933
transform 1 0 720 0 1 10101
box -29 -23 29 23
use L1M1_PR  L1M1_PR_399
timestamp 1626908933
transform 1 0 816 0 1 10175
box -29 -23 29 23
use L1M1_PR  L1M1_PR_297
timestamp 1626908933
transform 1 0 720 0 1 10101
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_136
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_424
timestamp 1626908933
transform 1 0 600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_284
timestamp 1626908933
transform 1 0 768 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_652
timestamp 1626908933
transform 1 0 768 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_12
timestamp 1626908933
transform 1 0 384 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_37
timestamp 1626908933
transform 1 0 384 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_0
timestamp 1626908933
transform 1 0 960 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_20
timestamp 1626908933
transform 1 0 960 0 -1 10656
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1093
timestamp 1626908933
transform 1 0 912 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_325
timestamp 1626908933
transform 1 0 912 0 1 10175
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1102
timestamp 1626908933
transform 1 0 1104 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_334
timestamp 1626908933
transform 1 0 1104 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_390
timestamp 1626908933
transform 1 0 1488 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1158
timestamp 1626908933
transform 1 0 1488 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_243
timestamp 1626908933
transform 1 0 1968 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1011
timestamp 1626908933
transform 1 0 1968 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_285
timestamp 1626908933
transform 1 0 1824 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_653
timestamp 1626908933
transform 1 0 1824 0 -1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_242
timestamp 1626908933
transform 1 0 1968 0 1 10101
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1010
timestamp 1626908933
transform 1 0 1968 0 1 10101
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_3
timestamp 1626908933
transform 1 0 1440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_12
timestamp 1626908933
transform 1 0 1440 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_41
timestamp 1626908933
transform 1 0 2016 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_16
timestamp 1626908933
transform 1 0 2016 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1142
timestamp 1626908933
transform 1 0 2400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_512
timestamp 1626908933
transform 1 0 2400 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_396
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_137
timestamp 1626908933
transform 1 0 2496 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_5
timestamp 1626908933
transform 1 0 2976 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_0
timestamp 1626908933
transform 1 0 2976 0 -1 10656
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1111
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_542
timestamp 1626908933
transform 1 0 2592 0 -1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_891
timestamp 1626908933
transform 1 0 3312 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_123
timestamp 1626908933
transform 1 0 3312 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1073
timestamp 1626908933
transform 1 0 3504 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_305
timestamp 1626908933
transform 1 0 3504 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1084
timestamp 1626908933
transform 1 0 3120 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_296
timestamp 1626908933
transform 1 0 3120 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_866
timestamp 1626908933
transform 1 0 3312 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_78
timestamp 1626908933
transform 1 0 3312 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1163
timestamp 1626908933
transform 1 0 3600 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_375
timestamp 1626908933
transform 1 0 3600 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1014
timestamp 1626908933
transform 1 0 3312 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_246
timestamp 1626908933
transform 1 0 3312 0 1 9805
box -32 -32 32 32
use M1M2_PR  M1M2_PR_831
timestamp 1626908933
transform 1 0 3504 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_63
timestamp 1626908933
transform 1 0 3504 0 1 9731
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_57
timestamp 1626908933
transform 1 0 3264 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_2
timestamp 1626908933
transform 1 0 3264 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1094
timestamp 1626908933
transform 1 0 3744 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_525
timestamp 1626908933
transform 1 0 3744 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_8
timestamp 1626908933
transform 1 0 4128 0 -1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_63
timestamp 1626908933
transform 1 0 4128 0 -1 10656
box -38 -49 518 715
use L1M1_PR  L1M1_PR_932
timestamp 1626908933
transform 1 0 3792 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_144
timestamp 1626908933
transform 1 0 3792 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_859
timestamp 1626908933
transform 1 0 4272 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_71
timestamp 1626908933
transform 1 0 4272 0 1 9657
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_382
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_112
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_382
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_112
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_382
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_112
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_120
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_408
timestamp 1626908933
transform 1 0 4600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_654
timestamp 1626908933
transform 1 0 4608 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_286
timestamp 1626908933
transform 1 0 4608 0 -1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_779
timestamp 1626908933
transform 1 0 4848 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1567
timestamp 1626908933
transform 1 0 4848 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_15
timestamp 1626908933
transform 1 0 4800 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_95
timestamp 1626908933
transform 1 0 4800 0 -1 10656
box -38 -49 902 715
use M1M2_PR  M1M2_PR_750
timestamp 1626908933
transform 1 0 5232 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1518
timestamp 1626908933
transform 1 0 5232 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_744
timestamp 1626908933
transform 1 0 6000 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1512
timestamp 1626908933
transform 1 0 6000 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_771
timestamp 1626908933
transform 1 0 6000 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1559
timestamp 1626908933
transform 1 0 6000 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_287
timestamp 1626908933
transform 1 0 5664 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_655
timestamp 1626908933
transform 1 0 5664 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_513
timestamp 1626908933
transform 1 0 5856 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1143
timestamp 1626908933
transform 1 0 5856 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_13
timestamp 1626908933
transform 1 0 5952 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_93
timestamp 1626908933
transform 1 0 5952 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_806
timestamp 1626908933
transform 1 0 6816 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_176
timestamp 1626908933
transform 1 0 6816 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1062
timestamp 1626908933
transform 1 0 6912 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_493
timestamp 1626908933
transform 1 0 6912 0 -1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_853
timestamp 1626908933
transform 1 0 6480 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_65
timestamp 1626908933
transform 1 0 6480 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_826
timestamp 1626908933
transform 1 0 6480 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_58
timestamp 1626908933
transform 1 0 6480 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_175
timestamp 1626908933
transform 1 0 7296 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_514
timestamp 1626908933
transform 1 0 7392 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_805
timestamp 1626908933
transform 1 0 7296 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1144
timestamp 1626908933
transform 1 0 7392 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_687
timestamp 1626908933
transform 1 0 7632 0 1 9583
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1455
timestamp 1626908933
transform 1 0 7632 0 1 9583
box -32 -32 32 32
use L1M1_PR  L1M1_PR_720
timestamp 1626908933
transform 1 0 7824 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1508
timestamp 1626908933
transform 1 0 7824 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_136
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_395
timestamp 1626908933
transform 1 0 7488 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_485
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1054
timestamp 1626908933
transform 1 0 7584 0 -1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_705
timestamp 1626908933
transform 1 0 7920 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1473
timestamp 1626908933
transform 1 0 7920 0 1 9509
box -32 -32 32 32
use M1M2_PR  M1M2_PR_114
timestamp 1626908933
transform 1 0 8112 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_882
timestamp 1626908933
transform 1 0 8112 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_133
timestamp 1626908933
transform 1 0 8112 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_921
timestamp 1626908933
transform 1 0 8112 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_515
timestamp 1626908933
transform 1 0 7968 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1145
timestamp 1626908933
transform 1 0 7968 0 -1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1523
timestamp 1626908933
transform 1 0 8688 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_735
timestamp 1626908933
transform 1 0 8688 0 1 9657
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_367
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_97
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_367
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_97
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_367
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_97
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_104
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_392
timestamp 1626908933
transform 1 0 8600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_10
timestamp 1626908933
transform 1 0 8064 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_90
timestamp 1626908933
transform 1 0 8064 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1046
timestamp 1626908933
transform 1 0 8928 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_476
timestamp 1626908933
transform 1 0 8928 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_87
timestamp 1626908933
transform 1 0 9696 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_7
timestamp 1626908933
transform 1 0 9696 0 -1 10656
box -38 -49 902 715
use L1M1_PR  L1M1_PR_915
timestamp 1626908933
transform 1 0 9072 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_127
timestamp 1626908933
transform 1 0 9072 0 1 9657
box -29 -23 29 23
use M1M2_PR  M1M2_PR_876
timestamp 1626908933
transform 1 0 9072 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_108
timestamp 1626908933
transform 1 0 9072 0 1 9657
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_804
timestamp 1626908933
transform 1 0 10560 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_174
timestamp 1626908933
transform 1 0 10560 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1453
timestamp 1626908933
transform 1 0 10320 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_685
timestamp 1626908933
transform 1 0 10320 0 1 9731
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_439
timestamp 1626908933
transform 1 0 10656 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1008
timestamp 1626908933
transform 1 0 10656 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_173
timestamp 1626908933
transform 1 0 11040 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_803
timestamp 1626908933
transform 1 0 11040 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_693
timestamp 1626908933
transform 1 0 11376 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1461
timestamp 1626908933
transform 1 0 11376 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_725
timestamp 1626908933
transform 1 0 11376 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1513
timestamp 1626908933
transform 1 0 11376 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_5
timestamp 1626908933
transform 1 0 11136 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_85
timestamp 1626908933
transform 1 0 11136 0 -1 10656
box -38 -49 902 715
use M1M2_PR  M1M2_PR_51
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -32 -32 32 32
use M1M2_PR  M1M2_PR_819
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -32 -32 32 32
use L1M1_PR  L1M1_PR_57
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -29 -23 29 23
use L1M1_PR  L1M1_PR_845
timestamp 1626908933
transform 1 0 11664 0 1 9657
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_172
timestamp 1626908933
transform 1 0 12000 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_802
timestamp 1626908933
transform 1 0 12000 0 -1 10656
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_352
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_82
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_352
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_82
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_352
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_82
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_376
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_88
timestamp 1626908933
transform 1 0 12600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_986
timestamp 1626908933
transform 1 0 12096 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_417
timestamp 1626908933
transform 1 0 12096 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_81
timestamp 1626908933
transform 1 0 12576 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_1
timestamp 1626908933
transform 1 0 12576 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_394
timestamp 1626908933
transform 1 0 12480 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_135
timestamp 1626908933
transform 1 0 12480 0 -1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1444
timestamp 1626908933
transform 1 0 13008 0 1 9731
box -32 -32 32 32
use M1M2_PR  M1M2_PR_676
timestamp 1626908933
transform 1 0 13008 0 1 9731
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_981
timestamp 1626908933
transform 1 0 14304 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_411
timestamp 1626908933
transform 1 0 14304 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_83
timestamp 1626908933
transform 1 0 13440 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_3
timestamp 1626908933
transform 1 0 13440 0 -1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_801
timestamp 1626908933
transform 1 0 15072 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_171
timestamp 1626908933
transform 1 0 15072 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_922
timestamp 1626908933
transform 1 0 15168 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_353
timestamp 1626908933
transform 1 0 15168 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_960
timestamp 1626908933
transform 1 0 15552 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_390
timestamp 1626908933
transform 1 0 15552 0 -1 10656
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_72
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_360
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_67
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_337
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_67
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_337
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_67
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_337
timestamp 1626908933
transform 1 0 16600 0 1 9990
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_328
timestamp 1626908933
transform 1 0 16320 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_897
timestamp 1626908933
transform 1 0 16320 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_364
timestamp 1626908933
transform 1 0 16704 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_934
timestamp 1626908933
transform 1 0 16704 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_393
timestamp 1626908933
transform 1 0 17472 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_134
timestamp 1626908933
transform 1 0 17472 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_872
timestamp 1626908933
transform 1 0 17760 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_303
timestamp 1626908933
transform 1 0 17760 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_478
timestamp 1626908933
transform 1 0 17568 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_110
timestamp 1626908933
transform 1 0 17568 0 -1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1384
timestamp 1626908933
transform 1 0 17232 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_616
timestamp 1626908933
transform 1 0 17232 0 1 9879
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_911
timestamp 1626908933
transform 1 0 18144 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_341
timestamp 1626908933
transform 1 0 18144 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_854
timestamp 1626908933
transform 1 0 18912 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_285
timestamp 1626908933
transform 1 0 18912 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_800
timestamp 1626908933
transform 1 0 19296 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_170
timestamp 1626908933
transform 1 0 19296 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_889
timestamp 1626908933
transform 1 0 19392 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_319
timestamp 1626908933
transform 1 0 19392 0 -1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_613
timestamp 1626908933
transform 1 0 19728 0 1 9879
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1381
timestamp 1626908933
transform 1 0 19728 0 1 9879
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_322
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_52
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_322
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_52
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_322
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_52
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_344
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_56
timestamp 1626908933
transform 1 0 20600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_477
timestamp 1626908933
transform 1 0 20160 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_109
timestamp 1626908933
transform 1 0 20160 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_269
timestamp 1626908933
transform 1 0 20352 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_838
timestamp 1626908933
transform 1 0 20352 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_860
timestamp 1626908933
transform 1 0 20736 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_290
timestamp 1626908933
transform 1 0 20736 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_476
timestamp 1626908933
transform 1 0 21504 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_108
timestamp 1626908933
transform 1 0 21504 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_836
timestamp 1626908933
transform 1 0 21696 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_266
timestamp 1626908933
transform 1 0 21696 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_819
timestamp 1626908933
transform 1 0 22656 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_249
timestamp 1626908933
transform 1 0 22656 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_799
timestamp 1626908933
transform 1 0 22560 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_169
timestamp 1626908933
transform 1 0 22560 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_392
timestamp 1626908933
transform 1 0 22464 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_133
timestamp 1626908933
transform 1 0 22464 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_796
timestamp 1626908933
transform 1 0 23424 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_226
timestamp 1626908933
transform 1 0 23424 0 -1 10656
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_307
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_37
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_307
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_37
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_307
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_37
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_328
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_40
timestamp 1626908933
transform 1 0 24600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_26
timestamp 1626908933
transform 1 0 25824 0 -1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_10
timestamp 1626908933
transform 1 0 25824 0 -1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_30
timestamp 1626908933
transform 1 0 24192 0 -1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_14
timestamp 1626908933
transform 1 0 24192 0 -1 10656
box -38 -49 1670 715
use M2M3_PR  M2M3_PR_105
timestamp 1626908933
transform 1 0 28080 0 1 9797
box -33 -37 33 37
use M2M3_PR  M2M3_PR_46
timestamp 1626908933
transform 1 0 28080 0 1 9797
box -33 -37 33 37
use osc_core_VIA7  osc_core_VIA7_292
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_22
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_292
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_22
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_292
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_22
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_312
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_24
timestamp 1626908933
transform 1 0 28600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_21
timestamp 1626908933
transform 1 0 27456 0 -1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_5
timestamp 1626908933
transform 1 0 27456 0 -1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_699
timestamp 1626908933
transform 1 0 29568 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_129
timestamp 1626908933
transform 1 0 29568 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_702
timestamp 1626908933
transform 1 0 29184 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_133
timestamp 1626908933
transform 1 0 29184 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_391
timestamp 1626908933
transform 1 0 29088 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_132
timestamp 1626908933
transform 1 0 29088 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_684
timestamp 1626908933
transform 1 0 30528 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_115
timestamp 1626908933
transform 1 0 30528 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_798
timestamp 1626908933
transform 1 0 30432 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_168
timestamp 1626908933
transform 1 0 30432 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_390
timestamp 1626908933
transform 1 0 30336 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_131
timestamp 1626908933
transform 1 0 30336 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_797
timestamp 1626908933
transform 1 0 30912 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_167
timestamp 1626908933
transform 1 0 30912 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_674
timestamp 1626908933
transform 1 0 31008 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_104
timestamp 1626908933
transform 1 0 31008 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_475
timestamp 1626908933
transform 1 0 31776 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_107
timestamp 1626908933
transform 1 0 31776 0 -1 10656
box -38 -49 230 715
use osc_core_VIA7  osc_core_VIA7_277
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_7
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_277
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_7
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_277
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_7
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_296
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_8
timestamp 1626908933
transform 1 0 32600 0 1 9990
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1146
timestamp 1626908933
transform 1 0 32352 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_516
timestamp 1626908933
transform 1 0 32352 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_389
timestamp 1626908933
transform 1 0 32448 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_130
timestamp 1626908933
transform 1 0 32448 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_65
timestamp 1626908933
transform 1 0 32544 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_634
timestamp 1626908933
transform 1 0 32544 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_82
timestamp 1626908933
transform 1 0 31968 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_651
timestamp 1626908933
transform 1 0 31968 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_629
timestamp 1626908933
transform 1 0 32928 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_59
timestamp 1626908933
transform 1 0 32928 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_796
timestamp 1626908933
transform 1 0 33696 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_166
timestamp 1626908933
transform 1 0 33696 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_601
timestamp 1626908933
transform 1 0 33792 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_32
timestamp 1626908933
transform 1 0 33792 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_599
timestamp 1626908933
transform 1 0 34176 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_29
timestamp 1626908933
transform 1 0 34176 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_7
timestamp 1626908933
transform 1 0 34944 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_577
timestamp 1626908933
transform 1 0 34944 0 -1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_662
timestamp 1626908933
transform 1 0 48 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_663
timestamp 1626908933
transform 1 0 240 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1430
timestamp 1626908933
transform 1 0 48 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1431
timestamp 1626908933
transform 1 0 240 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_659
timestamp 1626908933
transform 1 0 48 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1427
timestamp 1626908933
transform 1 0 48 0 1 10915
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_129
timestamp 1626908933
transform 1 0 288 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_388
timestamp 1626908933
transform 1 0 288 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_694
timestamp 1626908933
transform 1 0 432 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1482
timestamp 1626908933
transform 1 0 432 0 1 10397
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_288
timestamp 1626908933
transform 1 0 384 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_656
timestamp 1626908933
transform 1 0 384 0 1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1253
timestamp 1626908933
transform 1 0 816 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_465
timestamp 1626908933
transform 1 0 816 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1263
timestamp 1626908933
transform 1 0 528 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_475
timestamp 1626908933
transform 1 0 528 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1147
timestamp 1626908933
transform 1 0 576 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_517
timestamp 1626908933
transform 1 0 576 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_35
timestamp 1626908933
transform 1 0 672 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_10
timestamp 1626908933
transform 1 0 672 0 1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1252
timestamp 1626908933
transform 1 0 1104 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_464
timestamp 1626908933
transform 1 0 1104 0 1 10249
box -29 -23 29 23
use M2M3_PR  M2M3_PR_106
timestamp 1626908933
transform 1 0 1200 0 1 10285
box -33 -37 33 37
use M2M3_PR  M2M3_PR_47
timestamp 1626908933
transform 1 0 1200 0 1 10285
box -33 -37 33 37
use L1M1_PR  L1M1_PR_1461
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_673
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1409
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_641
timestamp 1626908933
transform 1 0 1200 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1248
timestamp 1626908933
transform 1 0 1392 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_460
timestamp 1626908933
transform 1 0 1392 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1195
timestamp 1626908933
transform 1 0 1008 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_407
timestamp 1626908933
transform 1 0 1008 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1103
timestamp 1626908933
transform 1 0 1008 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_335
timestamp 1626908933
transform 1 0 1008 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1479
timestamp 1626908933
transform 1 0 1104 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_691
timestamp 1626908933
transform 1 0 1104 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1105
timestamp 1626908933
transform 1 0 1296 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_337
timestamp 1626908933
transform 1 0 1296 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1200
timestamp 1626908933
transform 1 0 1392 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_412
timestamp 1626908933
transform 1 0 1392 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1249
timestamp 1626908933
transform 1 0 1200 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_461
timestamp 1626908933
transform 1 0 1200 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_11
timestamp 1626908933
transform 1 0 1056 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_36
timestamp 1626908933
transform 1 0 1056 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_625
timestamp 1626908933
transform 1 0 1440 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1255
timestamp 1626908933
transform 1 0 1440 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_1
timestamp 1626908933
transform 1 0 1536 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_0
timestamp 1626908933
transform 1 0 1536 0 1 10656
box -38 -49 230 715
use M1M2_PR  M1M2_PR_389
timestamp 1626908933
transform 1 0 1488 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1157
timestamp 1626908933
transform 1 0 1488 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_388
timestamp 1626908933
transform 1 0 1488 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1156
timestamp 1626908933
transform 1 0 1488 0 1 10989
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_550
timestamp 1626908933
transform 1 0 1728 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1119
timestamp 1626908933
transform 1 0 1728 0 1 10656
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1243
timestamp 1626908933
transform 1 0 2160 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_455
timestamp 1626908933
transform 1 0 2160 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1121
timestamp 1626908933
transform 1 0 2064 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_353
timestamp 1626908933
transform 1 0 2064 0 1 10397
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1214
timestamp 1626908933
transform 1 0 2352 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_426
timestamp 1626908933
transform 1 0 2352 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1098
timestamp 1626908933
transform 1 0 2352 0 1 10249
box -29 -23 29 23
use L1M1_PR  L1M1_PR_310
timestamp 1626908933
transform 1 0 2352 0 1 10249
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1429
timestamp 1626908933
transform 1 0 2160 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_661
timestamp 1626908933
transform 1 0 2160 0 1 10471
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1481
timestamp 1626908933
transform 1 0 1968 0 1 10471
box -29 -23 29 23
use L1M1_PR  L1M1_PR_693
timestamp 1626908933
transform 1 0 1968 0 1 10471
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_567
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_279
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_532
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_262
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_532
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_262
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_532
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_262
timestamp 1626908933
transform 1 0 2600 0 1 10656
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1083
timestamp 1626908933
transform 1 0 2352 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_295
timestamp 1626908933
transform 1 0 2352 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1207
timestamp 1626908933
transform 1 0 2448 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_419
timestamp 1626908933
transform 1 0 2448 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1112
timestamp 1626908933
transform 1 0 2352 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_344
timestamp 1626908933
transform 1 0 2352 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1480
timestamp 1626908933
transform 1 0 2160 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_692
timestamp 1626908933
transform 1 0 2160 0 1 10915
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1428
timestamp 1626908933
transform 1 0 2160 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_660
timestamp 1626908933
transform 1 0 2160 0 1 10915
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1241
timestamp 1626908933
transform 1 0 2256 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_453
timestamp 1626908933
transform 1 0 2256 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_165
timestamp 1626908933
transform 1 0 2496 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_795
timestamp 1626908933
transform 1 0 2496 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_15
timestamp 1626908933
transform 1 0 2112 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_40
timestamp 1626908933
transform 1 0 2112 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_1
timestamp 1626908933
transform 1 0 2976 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_56
timestamp 1626908933
transform 1 0 2976 0 1 10656
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1082
timestamp 1626908933
transform 1 0 3024 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_294
timestamp 1626908933
transform 1 0 3024 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1118
timestamp 1626908933
transform 1 0 2832 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_350
timestamp 1626908933
transform 1 0 2832 0 1 10397
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1110
timestamp 1626908933
transform 1 0 2592 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_541
timestamp 1626908933
transform 1 0 2592 0 1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1013
timestamp 1626908933
transform 1 0 3312 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_245
timestamp 1626908933
transform 1 0 3312 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1086
timestamp 1626908933
transform 1 0 3408 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_298
timestamp 1626908933
transform 1 0 3408 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_862
timestamp 1626908933
transform 1 0 3600 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_74
timestamp 1626908933
transform 1 0 3600 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1009
timestamp 1626908933
transform 1 0 3120 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_241
timestamp 1626908933
transform 1 0 3120 0 1 10397
box -32 -32 32 32
use L1M1_PR  L1M1_PR_867
timestamp 1626908933
transform 1 0 3216 0 1 10397
box -29 -23 29 23
use L1M1_PR  L1M1_PR_79
timestamp 1626908933
transform 1 0 3216 0 1 10397
box -29 -23 29 23
use M1M2_PR  M1M2_PR_830
timestamp 1626908933
transform 1 0 3504 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_62
timestamp 1626908933
transform 1 0 3504 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1008
timestamp 1626908933
transform 1 0 3120 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_240
timestamp 1626908933
transform 1 0 3120 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1012
timestamp 1626908933
transform 1 0 3312 0 1 10841
box -32 -32 32 32
use M1M2_PR  M1M2_PR_244
timestamp 1626908933
transform 1 0 3312 0 1 10841
box -32 -32 32 32
use M1M2_PR  M1M2_PR_834
timestamp 1626908933
transform 1 0 3312 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_66
timestamp 1626908933
transform 1 0 3312 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1087
timestamp 1626908933
transform 1 0 3216 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_865
timestamp 1626908933
transform 1 0 3312 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_299
timestamp 1626908933
transform 1 0 3216 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_77
timestamp 1626908933
transform 1 0 3312 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_829
timestamp 1626908933
transform 1 0 3504 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_61
timestamp 1626908933
transform 1 0 3504 0 1 10915
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_58
timestamp 1626908933
transform 1 0 3456 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_3
timestamp 1626908933
transform 1 0 3456 0 1 10656
box -38 -49 518 715
use M1M2_PR  M1M2_PR_247
timestamp 1626908933
transform 1 0 3696 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1015
timestamp 1626908933
transform 1 0 3696 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_73
timestamp 1626908933
transform 1 0 3792 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_301
timestamp 1626908933
transform 1 0 3696 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_861
timestamp 1626908933
transform 1 0 3792 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1089
timestamp 1626908933
transform 1 0 3696 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_518
timestamp 1626908933
transform 1 0 3936 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1148
timestamp 1626908933
transform 1 0 3936 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_62
timestamp 1626908933
transform 1 0 4032 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_7
timestamp 1626908933
transform 1 0 4032 0 1 10656
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1097
timestamp 1626908933
transform 1 0 4272 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_309
timestamp 1626908933
transform 1 0 4272 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_857
timestamp 1626908933
transform 1 0 4464 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_69
timestamp 1626908933
transform 1 0 4464 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1021
timestamp 1626908933
transform 1 0 4368 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_253
timestamp 1626908933
transform 1 0 4368 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1096
timestamp 1626908933
transform 1 0 4272 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_308
timestamp 1626908933
transform 1 0 4272 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_858
timestamp 1626908933
transform 1 0 4368 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_70
timestamp 1626908933
transform 1 0 4368 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_128
timestamp 1626908933
transform 1 0 4992 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_387
timestamp 1626908933
transform 1 0 4992 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_306
timestamp 1626908933
transform 1 0 4656 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1094
timestamp 1626908933
transform 1 0 4656 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_59
timestamp 1626908933
transform 1 0 4848 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_827
timestamp 1626908933
transform 1 0 4848 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_67
timestamp 1626908933
transform 1 0 4848 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_855
timestamp 1626908933
transform 1 0 4848 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_65
timestamp 1626908933
transform 1 0 4512 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_10
timestamp 1626908933
transform 1 0 4512 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_164
timestamp 1626908933
transform 1 0 5088 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_794
timestamp 1626908933
transform 1 0 5088 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_749
timestamp 1626908933
transform 1 0 5232 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1517
timestamp 1626908933
transform 1 0 5232 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_66
timestamp 1626908933
transform 1 0 5328 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_776
timestamp 1626908933
transform 1 0 5232 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_854
timestamp 1626908933
transform 1 0 5328 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1564
timestamp 1626908933
transform 1 0 5232 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_520
timestamp 1626908933
transform 1 0 5184 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1090
timestamp 1626908933
transform 1 0 5184 0 1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1511
timestamp 1626908933
transform 1 0 6000 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_743
timestamp 1626908933
transform 1 0 6000 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1556
timestamp 1626908933
transform 1 0 6096 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_768
timestamp 1626908933
transform 1 0 6096 0 1 10323
box -29 -23 29 23
use M2M3_PR  M2M3_PR_117
timestamp 1626908933
transform 1 0 6000 0 1 10895
box -33 -37 33 37
use M2M3_PR  M2M3_PR_58
timestamp 1626908933
transform 1 0 6000 0 1 10895
box -33 -37 33 37
use L1M1_PR  L1M1_PR_1104
timestamp 1626908933
transform 1 0 6096 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_316
timestamp 1626908933
transform 1 0 6096 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1026
timestamp 1626908933
transform 1 0 6096 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_258
timestamp 1626908933
transform 1 0 6096 0 1 10989
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_263
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_551
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -142 200 178
use L1M1_PR  L1M1_PR_852
timestamp 1626908933
transform 1 0 6480 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_64
timestamp 1626908933
transform 1 0 6480 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_825
timestamp 1626908933
transform 1 0 6480 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_57
timestamp 1626908933
transform 1 0 6480 0 1 10323
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_247
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_517
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_247
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_517
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_247
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_517
timestamp 1626908933
transform 1 0 6600 0 1 10656
box -200 -49 200 49
use M1M2_PR  M1M2_PR_29
timestamp 1626908933
transform 1 0 6384 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_797
timestamp 1626908933
transform 1 0 6384 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_36
timestamp 1626908933
transform 1 0 6288 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_824
timestamp 1626908933
transform 1 0 6288 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_793
timestamp 1626908933
transform 1 0 6432 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_163
timestamp 1626908933
transform 1 0 6432 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_496
timestamp 1626908933
transform 1 0 6528 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1065
timestamp 1626908933
transform 1 0 6528 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_67
timestamp 1626908933
transform 1 0 5952 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_12
timestamp 1626908933
transform 1 0 5952 0 1 10656
box -38 -49 518 715
use M2M3_PR  M2M3_PR_116
timestamp 1626908933
transform 1 0 6864 0 1 10895
box -33 -37 33 37
use M2M3_PR  M2M3_PR_57
timestamp 1626908933
transform 1 0 6864 0 1 10895
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_792
timestamp 1626908933
transform 1 0 6912 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_162
timestamp 1626908933
transform 1 0 6912 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_56
timestamp 1626908933
transform 1 0 7056 0 1 10397
box -32 -32 32 32
use M1M2_PR  M1M2_PR_824
timestamp 1626908933
transform 1 0 7056 0 1 10397
box -32 -32 32 32
use L1M1_PR  L1M1_PR_758
timestamp 1626908933
transform 1 0 7728 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1546
timestamp 1626908933
transform 1 0 7728 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_55
timestamp 1626908933
transform 1 0 7056 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_823
timestamp 1626908933
transform 1 0 7056 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_63
timestamp 1626908933
transform 1 0 7152 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_851
timestamp 1626908933
transform 1 0 7152 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_489
timestamp 1626908933
transform 1 0 7872 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1059
timestamp 1626908933
transform 1 0 7872 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_9
timestamp 1626908933
transform -1 0 7872 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_89
timestamp 1626908933
transform -1 0 7872 0 1 10656
box -38 -49 902 715
use M1M2_PR  M1M2_PR_727
timestamp 1626908933
transform 1 0 8304 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1495
timestamp 1626908933
transform 1 0 8304 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_756
timestamp 1626908933
transform 1 0 8304 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1544
timestamp 1626908933
transform 1 0 8304 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_726
timestamp 1626908933
transform 1 0 8304 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1494
timestamp 1626908933
transform 1 0 8304 0 1 10989
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_289
timestamp 1626908933
transform 1 0 8640 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_657
timestamp 1626908933
transform 1 0 8640 0 1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_62
timestamp 1626908933
transform 1 0 8592 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_850
timestamp 1626908933
transform 1 0 8592 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_519
timestamp 1626908933
transform 1 0 8832 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1149
timestamp 1626908933
transform 1 0 8832 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_54
timestamp 1626908933
transform 1 0 8880 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_822
timestamp 1626908933
transform 1 0 8880 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_52
timestamp 1626908933
transform 1 0 9168 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_820
timestamp 1626908933
transform 1 0 9168 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_750
timestamp 1626908933
transform 1 0 9072 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1538
timestamp 1626908933
transform 1 0 9072 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_60
timestamp 1626908933
transform 1 0 9648 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_848
timestamp 1626908933
transform 1 0 9648 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_8
timestamp 1626908933
transform 1 0 8928 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_88
timestamp 1626908933
transform 1 0 8928 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_127
timestamp 1626908933
transform 1 0 9984 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_386
timestamp 1626908933
transform 1 0 9984 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_290
timestamp 1626908933
transform 1 0 9792 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_658
timestamp 1626908933
transform 1 0 9792 0 1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_732
timestamp 1626908933
transform 1 0 9936 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1520
timestamp 1626908933
transform 1 0 9936 0 1 10323
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_247
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_535
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -142 200 178
use L1M1_PR  L1M1_PR_847
timestamp 1626908933
transform 1 0 10224 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_59
timestamp 1626908933
transform 1 0 10224 0 1 10323
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_502
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_232
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_502
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_232
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_502
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_232
timestamp 1626908933
transform 1 0 10600 0 1 10656
box -200 -49 200 49
use L1M1_PR  L1M1_PR_846
timestamp 1626908933
transform 1 0 10224 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_58
timestamp 1626908933
transform 1 0 10224 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_6
timestamp 1626908933
transform -1 0 10944 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_86
timestamp 1626908933
transform -1 0 10944 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_161
timestamp 1626908933
transform 1 0 10944 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_791
timestamp 1626908933
transform 1 0 10944 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_699
timestamp 1626908933
transform 1 0 10992 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1467
timestamp 1626908933
transform 1 0 10992 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_698
timestamp 1626908933
transform 1 0 10992 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1466
timestamp 1626908933
transform 1 0 10992 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_730
timestamp 1626908933
transform 1 0 10800 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1518
timestamp 1626908933
transform 1 0 10800 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_692
timestamp 1626908933
transform 1 0 11376 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1460
timestamp 1626908933
transform 1 0 11376 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_726
timestamp 1626908933
transform 1 0 11280 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1514
timestamp 1626908933
transform 1 0 11280 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_454
timestamp 1626908933
transform 1 0 11040 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1024
timestamp 1626908933
transform 1 0 11040 0 1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_50
timestamp 1626908933
transform 1 0 11664 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_818
timestamp 1626908933
transform 1 0 11664 0 1 10323
box -32 -32 32 32
use L1M1_PR  L1M1_PR_56
timestamp 1626908933
transform 1 0 11664 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_844
timestamp 1626908933
transform 1 0 11664 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_21
timestamp 1626908933
transform 1 0 12336 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_789
timestamp 1626908933
transform 1 0 12336 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_15
timestamp 1626908933
transform 1 0 12336 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_803
timestamp 1626908933
transform 1 0 12336 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_722
timestamp 1626908933
transform 1 0 11952 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1510
timestamp 1626908933
transform 1 0 11952 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_20
timestamp 1626908933
transform 1 0 11808 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_100
timestamp 1626908933
transform 1 0 11808 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_291
timestamp 1626908933
transform 1 0 12672 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_659
timestamp 1626908933
transform 1 0 12672 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_520
timestamp 1626908933
transform 1 0 12864 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1150
timestamp 1626908933
transform 1 0 12864 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_708
timestamp 1626908933
transform 1 0 12816 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1496
timestamp 1626908933
transform 1 0 12816 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_675
timestamp 1626908933
transform 1 0 13008 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1443
timestamp 1626908933
transform 1 0 13008 0 1 10249
box -32 -32 32 32
use L1M1_PR  L1M1_PR_55
timestamp 1626908933
transform 1 0 13104 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_843
timestamp 1626908933
transform 1 0 13104 0 1 10323
box -29 -23 29 23
use M1M2_PR  M1M2_PR_674
timestamp 1626908933
transform 1 0 13104 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1442
timestamp 1626908933
transform 1 0 13104 0 1 10989
box -32 -32 32 32
use L1M1_PR  L1M1_PR_707
timestamp 1626908933
transform 1 0 13104 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1495
timestamp 1626908933
transform 1 0 13104 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_2
timestamp 1626908933
transform 1 0 12960 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_82
timestamp 1626908933
transform 1 0 12960 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_292
timestamp 1626908933
transform 1 0 13824 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_660
timestamp 1626908933
transform 1 0 13824 0 1 10656
box -38 -49 230 715
use L1M1_PR  L1M1_PR_705
timestamp 1626908933
transform 1 0 13584 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1493
timestamp 1626908933
transform 1 0 13584 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_54
timestamp 1626908933
transform 1 0 13680 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_842
timestamp 1626908933
transform 1 0 13680 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_841
timestamp 1626908933
transform 1 0 13968 0 1 10323
box -29 -23 29 23
use L1M1_PR  L1M1_PR_53
timestamp 1626908933
transform 1 0 13968 0 1 10323
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1151
timestamp 1626908933
transform 1 0 14016 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_521
timestamp 1626908933
transform 1 0 14016 0 1 10656
box -38 -49 134 715
use M2M3_PR_R  M2M3_PR_R_2
timestamp 1626908933
transform 1 0 14064 0 1 10895
box -37 -33 37 33
use M2M3_PR_R  M2M3_PR_R_0
timestamp 1626908933
transform 1 0 14064 0 1 10895
box -37 -33 37 33
use M1M2_PR  M1M2_PR_816
timestamp 1626908933
transform 1 0 14064 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_48
timestamp 1626908933
transform 1 0 14064 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_817
timestamp 1626908933
transform 1 0 14064 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_49
timestamp 1626908933
transform 1 0 14064 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_0
timestamp 1626908933
transform 1 0 14112 0 1 10656
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_80
timestamp 1626908933
transform 1 0 14112 0 1 10656
box -38 -49 902 715
use osc_core_VIA4  osc_core_VIA4_231
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_519
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_487
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_217
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_487
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_217
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_487
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_217
timestamp 1626908933
transform 1 0 14600 0 1 10656
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1491
timestamp 1626908933
transform 1 0 14352 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_840
timestamp 1626908933
transform 1 0 14640 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_703
timestamp 1626908933
transform 1 0 14352 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_52
timestamp 1626908933
transform 1 0 14640 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_352
timestamp 1626908933
transform 1 0 15168 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_921
timestamp 1626908933
transform 1 0 15168 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_160
timestamp 1626908933
transform 1 0 15072 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_790
timestamp 1626908933
transform 1 0 15072 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_126
timestamp 1626908933
transform 1 0 14976 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_385
timestamp 1626908933
transform 1 0 14976 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_959
timestamp 1626908933
transform 1 0 15552 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_389
timestamp 1626908933
transform 1 0 15552 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_933
timestamp 1626908933
transform 1 0 16896 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_363
timestamp 1626908933
transform 1 0 16896 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_474
timestamp 1626908933
transform 1 0 16320 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_106
timestamp 1626908933
transform 1 0 16320 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_896
timestamp 1626908933
transform 1 0 16512 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_327
timestamp 1626908933
transform 1 0 16512 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_871
timestamp 1626908933
transform 1 0 17760 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_302
timestamp 1626908933
transform 1 0 17760 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_789
timestamp 1626908933
transform 1 0 17664 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_159
timestamp 1626908933
transform 1 0 17664 0 1 10656
box -38 -49 134 715
use M3M4_PR  M3M4_PR_25
timestamp 1626908933
transform 1 0 17904 0 1 10895
box -38 -33 38 33
use M3M4_PR  M3M4_PR_4
timestamp 1626908933
transform 1 0 17904 0 1 10895
box -38 -33 38 33
use M1M2_PR  M1M2_PR_1324
timestamp 1626908933
transform 1 0 17904 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_556
timestamp 1626908933
transform 1 0 17904 0 1 10249
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_503
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_215
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_202
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_472
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_202
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_472
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_202
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_472
timestamp 1626908933
transform 1 0 18600 0 1 10656
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_340
timestamp 1626908933
transform 1 0 18144 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_910
timestamp 1626908933
transform 1 0 18144 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_788
timestamp 1626908933
transform 1 0 19104 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_158
timestamp 1626908933
transform 1 0 19104 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_473
timestamp 1626908933
transform 1 0 18912 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_105
timestamp 1626908933
transform 1 0 18912 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_888
timestamp 1626908933
transform 1 0 19200 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_318
timestamp 1626908933
transform 1 0 19200 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_871
timestamp 1626908933
transform 1 0 20064 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_301
timestamp 1626908933
transform 1 0 20064 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_384
timestamp 1626908933
transform 1 0 19968 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_125
timestamp 1626908933
transform 1 0 19968 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_822
timestamp 1626908933
transform 1 0 21024 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_253
timestamp 1626908933
transform 1 0 21024 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_472
timestamp 1626908933
transform 1 0 20832 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_104
timestamp 1626908933
transform 1 0 20832 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_845
timestamp 1626908933
transform 1 0 21408 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_275
timestamp 1626908933
transform 1 0 21408 0 1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_555
timestamp 1626908933
transform 1 0 21936 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1323
timestamp 1626908933
transform 1 0 21936 0 1 10249
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_199
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_487
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_187
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_457
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_187
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_457
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_187
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_457
timestamp 1626908933
transform 1 0 22600 0 1 10656
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_234
timestamp 1626908933
transform 1 0 22176 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_803
timestamp 1626908933
transform 1 0 22176 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_818
timestamp 1626908933
transform 1 0 22560 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_248
timestamp 1626908933
transform 1 0 22560 0 1 10656
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1342
timestamp 1626908933
transform 1 0 23472 0 1 10915
box -29 -23 29 23
use L1M1_PR  L1M1_PR_554
timestamp 1626908933
transform 1 0 23472 0 1 10915
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_63
timestamp 1626908933
transform 1 0 23328 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_23
timestamp 1626908933
transform 1 0 23328 0 1 10656
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1254
timestamp 1626908933
transform 1 0 23664 0 1 10915
box -32 -32 32 32
use M1M2_PR  M1M2_PR_486
timestamp 1626908933
transform 1 0 23664 0 1 10915
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_383
timestamp 1626908933
transform 1 0 24096 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_124
timestamp 1626908933
transform 1 0 24096 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1133
timestamp 1626908933
transform 1 0 23856 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_365
timestamp 1626908933
transform 1 0 23856 0 1 10249
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_29
timestamp 1626908933
transform 1 0 25824 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_9
timestamp 1626908933
transform 1 0 25824 0 1 10656
box -38 -49 518 715
use M1M2_PR  M1M2_PR_439
timestamp 1626908933
transform 1 0 25776 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1207
timestamp 1626908933
transform 1 0 25776 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_438
timestamp 1626908933
transform 1 0 25776 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1206
timestamp 1626908933
transform 1 0 25776 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1203
timestamp 1626908933
transform 1 0 26160 0 1 10471
box -32 -32 32 32
use M1M2_PR  M1M2_PR_435
timestamp 1626908933
transform 1 0 26160 0 1 10471
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1287
timestamp 1626908933
transform 1 0 26160 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_499
timestamp 1626908933
transform 1 0 26160 0 1 10767
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1202
timestamp 1626908933
transform 1 0 26160 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_434
timestamp 1626908933
transform 1 0 26160 0 1 10767
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1285
timestamp 1626908933
transform 1 0 26160 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_497
timestamp 1626908933
transform 1 0 26160 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1201
timestamp 1626908933
transform 1 0 26160 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_433
timestamp 1626908933
transform 1 0 26160 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1274
timestamp 1626908933
transform 1 0 26256 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_506
timestamp 1626908933
transform 1 0 26256 0 1 10989
box -32 -32 32 32
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_29
timestamp 1626908933
transform 1 0 24192 0 1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_13
timestamp 1626908933
transform 1 0 24192 0 1 10656
box -38 -49 1670 715
use osc_core_VIA4  osc_core_VIA4_183
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_471
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_442
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_172
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_442
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_172
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_442
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_172
timestamp 1626908933
transform 1 0 26600 0 1 10656
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1365
timestamp 1626908933
transform 1 0 26352 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_577
timestamp 1626908933
transform 1 0 26352 0 1 10989
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_293
timestamp 1626908933
transform 1 0 27072 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_661
timestamp 1626908933
transform 1 0 27072 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_39
timestamp 1626908933
transform 1 0 26304 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_79
timestamp 1626908933
transform 1 0 26304 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1152
timestamp 1626908933
transform 1 0 27264 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_522
timestamp 1626908933
transform 1 0 27264 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_382
timestamp 1626908933
transform 1 0 27360 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_123
timestamp 1626908933
transform 1 0 27360 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1278
timestamp 1626908933
transform 1 0 27504 0 1 10989
box -29 -23 29 23
use L1M1_PR  L1M1_PR_490
timestamp 1626908933
transform 1 0 27504 0 1 10989
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1188
timestamp 1626908933
transform 1 0 27504 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_420
timestamp 1626908933
transform 1 0 27504 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1189
timestamp 1626908933
transform 1 0 27504 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_421
timestamp 1626908933
transform 1 0 27504 0 1 10767
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1190
timestamp 1626908933
transform 1 0 27504 0 1 10323
box -32 -32 32 32
use M1M2_PR  M1M2_PR_422
timestamp 1626908933
transform 1 0 27504 0 1 10323
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_157
timestamp 1626908933
transform 1 0 27936 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_787
timestamp 1626908933
transform 1 0 27936 0 1 10656
box -38 -49 134 715
use L1M1_PR  L1M1_PR_491
timestamp 1626908933
transform 1 0 27600 0 1 10767
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1279
timestamp 1626908933
transform 1 0 27600 0 1 10767
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_28
timestamp 1626908933
transform 1 0 27456 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_8
timestamp 1626908933
transform 1 0 27456 0 1 10656
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_723
timestamp 1626908933
transform 1 0 28416 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_153
timestamp 1626908933
transform 1 0 28416 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_727
timestamp 1626908933
transform 1 0 28032 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_158
timestamp 1626908933
transform 1 0 28032 0 1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1195
timestamp 1626908933
transform 1 0 29040 0 1 10249
box -32 -32 32 32
use M1M2_PR  M1M2_PR_427
timestamp 1626908933
transform 1 0 29040 0 1 10249
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_132
timestamp 1626908933
transform 1 0 29184 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_701
timestamp 1626908933
transform 1 0 29184 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_122
timestamp 1626908933
transform 1 0 29568 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_381
timestamp 1626908933
transform 1 0 29568 0 1 10656
box -38 -49 134 715
use M1M2_PR  M1M2_PR_416
timestamp 1626908933
transform 1 0 29712 0 1 10989
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1184
timestamp 1626908933
transform 1 0 29712 0 1 10989
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_157
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_427
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_157
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_427
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_157
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_427
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_167
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_455
timestamp 1626908933
transform 1 0 30600 0 1 10656
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_666
timestamp 1626908933
transform 1 0 31296 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_97
timestamp 1626908933
transform 1 0 31296 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_658
timestamp 1626908933
transform 1 0 31680 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_88
timestamp 1626908933
transform 1 0 31680 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_20
timestamp 1626908933
transform 1 0 29664 0 1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_4
timestamp 1626908933
transform 1 0 29664 0 1 10656
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_633
timestamp 1626908933
transform 1 0 32544 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_64
timestamp 1626908933
transform 1 0 32544 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_786
timestamp 1626908933
transform 1 0 32448 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_156
timestamp 1626908933
transform 1 0 32448 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_628
timestamp 1626908933
transform 1 0 32928 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_58
timestamp 1626908933
transform 1 0 32928 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_785
timestamp 1626908933
transform 1 0 33696 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_155
timestamp 1626908933
transform 1 0 33696 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_600
timestamp 1626908933
transform 1 0 33792 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_31
timestamp 1626908933
transform 1 0 33792 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_598
timestamp 1626908933
transform 1 0 34176 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_28
timestamp 1626908933
transform 1 0 34176 0 1 10656
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_412
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_142
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_412
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_142
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_412
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_142
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_151
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_439
timestamp 1626908933
transform 1 0 34600 0 1 10656
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_121
timestamp 1626908933
transform 1 0 34944 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_380
timestamp 1626908933
transform 1 0 34944 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_294
timestamp 1626908933
transform 1 0 35424 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_662
timestamp 1626908933
transform 1 0 35424 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_523
timestamp 1626908933
transform 1 0 35616 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1153
timestamp 1626908933
transform 1 0 35616 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_7
timestamp 1626908933
transform 1 0 35040 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_576
timestamp 1626908933
transform 1 0 35040 0 1 10656
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1426
timestamp 1626908933
transform 1 0 144 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_658
timestamp 1626908933
transform 1 0 144 0 1 11211
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_396
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_126
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_396
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_126
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_396
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_126
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_423
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_135
timestamp 1626908933
transform 1 0 600 0 1 11322
box -200 -142 200 178
use M1M2_PR  M1M2_PR_657
timestamp 1626908933
transform 1 0 48 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1425
timestamp 1626908933
transform 1 0 48 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_689
timestamp 1626908933
transform 1 0 432 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1477
timestamp 1626908933
transform 1 0 432 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_524
timestamp 1626908933
transform 1 0 288 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1154
timestamp 1626908933
transform 1 0 288 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_9
timestamp 1626908933
transform 1 0 384 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_34
timestamp 1626908933
transform 1 0 384 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_690
timestamp 1626908933
transform 1 0 624 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1478
timestamp 1626908933
transform 1 0 624 0 1 11211
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1038
timestamp 1626908933
transform 1 0 624 0 1 11507
box -32 -32 32 32
use M1M2_PR  M1M2_PR_270
timestamp 1626908933
transform 1 0 624 0 1 11507
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1102
timestamp 1626908933
transform 1 0 720 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_314
timestamp 1626908933
transform 1 0 720 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1262
timestamp 1626908933
transform 1 0 528 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_474
timestamp 1626908933
transform 1 0 528 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1190
timestamp 1626908933
transform 1 0 720 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_402
timestamp 1626908933
transform 1 0 720 0 1 11729
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1097
timestamp 1626908933
transform 1 0 720 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_329
timestamp 1626908933
transform 1 0 720 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1160
timestamp 1626908933
transform 1 0 912 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_392
timestamp 1626908933
transform 1 0 912 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_295
timestamp 1626908933
transform 1 0 768 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_663
timestamp 1626908933
transform 1 0 768 0 -1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_317
timestamp 1626908933
transform 1 0 1008 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1105
timestamp 1626908933
transform 1 0 1008 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_463
timestamp 1626908933
transform 1 0 1104 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1251
timestamp 1626908933
transform 1 0 1104 0 1 11655
box -29 -23 29 23
use M2M3_PR  M2M3_PR_80
timestamp 1626908933
transform 1 0 1200 0 1 11139
box -33 -37 33 37
use M2M3_PR  M2M3_PR_21
timestamp 1626908933
transform 1 0 1200 0 1 11139
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1027
timestamp 1626908933
transform 1 0 1200 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_259
timestamp 1626908933
transform 1 0 1200 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1110
timestamp 1626908933
transform 1 0 1392 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_322
timestamp 1626908933
transform 1 0 1392 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1194
timestamp 1626908933
transform 1 0 1296 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_406
timestamp 1626908933
transform 1 0 1296 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1155
timestamp 1626908933
transform 1 0 1344 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_525
timestamp 1626908933
transform 1 0 1344 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_7
timestamp 1626908933
transform 1 0 960 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_32
timestamp 1626908933
transform 1 0 960 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1224
timestamp 1626908933
transform 1 0 1584 0 1 11137
box -32 -32 32 32
use M1M2_PR  M1M2_PR_456
timestamp 1626908933
transform 1 0 1584 0 1 11137
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1302
timestamp 1626908933
transform 1 0 1584 0 1 11137
box -29 -23 29 23
use L1M1_PR  L1M1_PR_514
timestamp 1626908933
transform 1 0 1584 0 1 11137
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1155
timestamp 1626908933
transform 1 0 1488 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_387
timestamp 1626908933
transform 1 0 1488 0 1 11655
box -32 -32 32 32
use M3M4_PR  M3M4_PR_40
timestamp 1626908933
transform 1 0 1632 0 1 11627
box -38 -33 38 33
use M3M4_PR  M3M4_PR_19
timestamp 1626908933
transform 1 0 1632 0 1 11627
box -38 -33 38 33
use M2M3_PR  M2M3_PR_87
timestamp 1626908933
transform 1 0 1584 0 1 11627
box -33 -37 33 37
use M2M3_PR  M2M3_PR_28
timestamp 1626908933
transform 1 0 1584 0 1 11627
box -33 -37 33 37
use L1M1_PR  L1M1_PR_1301
timestamp 1626908933
transform 1 0 1584 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_513
timestamp 1626908933
transform 1 0 1584 0 1 11729
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1223
timestamp 1626908933
transform 1 0 1584 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_455
timestamp 1626908933
transform 1 0 1584 0 1 11729
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_526
timestamp 1626908933
transform 1 0 2016 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1156
timestamp 1626908933
transform 1 0 2016 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_3
timestamp 1626908933
transform -1 0 2016 0 -1 11988
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_4  sky130_fd_sc_hs__clkbuf_4_0
timestamp 1626908933
transform -1 0 2016 0 -1 11988
box -38 -49 614 715
use M1M2_PR  M1M2_PR_343
timestamp 1626908933
transform 1 0 2352 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1111
timestamp 1626908933
transform 1 0 2352 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_452
timestamp 1626908933
transform 1 0 2256 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1240
timestamp 1626908933
transform 1 0 2256 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_120
timestamp 1626908933
transform 1 0 2496 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_379
timestamp 1626908933
transform 1 0 2496 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_418
timestamp 1626908933
transform 1 0 2448 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1206
timestamp 1626908933
transform 1 0 2448 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_77
timestamp 1626908933
transform 1 0 2592 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_22
timestamp 1626908933
transform 1 0 2592 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_17
timestamp 1626908933
transform 1 0 2112 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_42
timestamp 1626908933
transform 1 0 2112 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_330
timestamp 1626908933
transform 1 0 2736 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1118
timestamp 1626908933
transform 1 0 2736 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_96
timestamp 1626908933
transform 1 0 2928 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_864
timestamp 1626908933
transform 1 0 2928 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_112
timestamp 1626908933
transform 1 0 2928 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_900
timestamp 1626908933
transform 1 0 2928 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_527
timestamp 1626908933
transform 1 0 3072 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1157
timestamp 1626908933
transform 1 0 3072 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_65
timestamp 1626908933
transform 1 0 3312 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_833
timestamp 1626908933
transform 1 0 3312 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_76
timestamp 1626908933
transform 1 0 3312 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_864
timestamp 1626908933
transform 1 0 3312 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_60
timestamp 1626908933
transform -1 0 3648 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_5
timestamp 1626908933
transform -1 0 3648 0 -1 11988
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1091
timestamp 1626908933
transform 1 0 3504 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_303
timestamp 1626908933
transform 1 0 3504 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1018
timestamp 1626908933
transform 1 0 3504 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_250
timestamp 1626908933
transform 1 0 3504 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1093
timestamp 1626908933
transform 1 0 3840 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_524
timestamp 1626908933
transform 1 0 3840 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_471
timestamp 1626908933
transform 1 0 3648 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_103
timestamp 1626908933
transform 1 0 3648 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1020
timestamp 1626908933
transform 1 0 4464 0 1 11063
box -32 -32 32 32
use M1M2_PR  M1M2_PR_252
timestamp 1626908933
transform 1 0 4464 0 1 11063
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_381
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_111
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_381
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_111
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_381
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_111
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_119
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_407
timestamp 1626908933
transform 1 0 4600 0 1 11322
box -200 -142 200 178
use L1M1_PR  L1M1_PR_68
timestamp 1626908933
transform 1 0 4560 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_856
timestamp 1626908933
transform 1 0 4560 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_254
timestamp 1626908933
transform 1 0 4272 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1022
timestamp 1626908933
transform 1 0 4272 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_307
timestamp 1626908933
transform 1 0 4368 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1095
timestamp 1626908933
transform 1 0 4368 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_296
timestamp 1626908933
transform 1 0 4704 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_664
timestamp 1626908933
transform 1 0 4704 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_64
timestamp 1626908933
transform 1 0 4224 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_9
timestamp 1626908933
transform 1 0 4224 0 -1 11988
box -38 -49 518 715
use M1M2_PR  M1M2_PR_828
timestamp 1626908933
transform 1 0 4752 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_60
timestamp 1626908933
transform 1 0 4752 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1124
timestamp 1626908933
transform 1 0 5136 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_336
timestamp 1626908933
transform 1 0 5136 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_28
timestamp 1626908933
transform 1 0 4992 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_83
timestamp 1626908933
transform 1 0 4992 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1158
timestamp 1626908933
transform 1 0 4896 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_528
timestamp 1626908933
transform 1 0 4896 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_297
timestamp 1626908933
transform 1 0 5472 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_665
timestamp 1626908933
transform 1 0 5472 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_84
timestamp 1626908933
transform 1 0 5328 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_852
timestamp 1626908933
transform 1 0 5328 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_100
timestamp 1626908933
transform 1 0 5328 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_888
timestamp 1626908933
transform 1 0 5328 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_529
timestamp 1626908933
transform 1 0 5664 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1159
timestamp 1626908933
transform 1 0 5664 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_256
timestamp 1626908933
transform 1 0 5616 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1024
timestamp 1626908933
transform 1 0 5616 0 1 11581
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_1
timestamp 1626908933
transform 1 0 5760 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_6
timestamp 1626908933
transform 1 0 5760 0 -1 11988
box -38 -49 326 715
use M2M3_PR  M2M3_PR_20
timestamp 1626908933
transform 1 0 6096 0 1 11139
box -33 -37 33 37
use M2M3_PR  M2M3_PR_79
timestamp 1626908933
transform 1 0 6096 0 1 11139
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1025
timestamp 1626908933
transform 1 0 6096 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_257
timestamp 1626908933
transform 1 0 6096 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1103
timestamp 1626908933
transform 1 0 6192 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_315
timestamp 1626908933
transform 1 0 6192 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_821
timestamp 1626908933
transform 1 0 6384 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_33
timestamp 1626908933
transform 1 0 6384 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_796
timestamp 1626908933
transform 1 0 6384 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_28
timestamp 1626908933
transform 1 0 6384 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_827
timestamp 1626908933
transform 1 0 6000 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_39
timestamp 1626908933
transform 1 0 6000 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_68
timestamp 1626908933
transform 1 0 6048 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_13
timestamp 1626908933
transform 1 0 6048 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1064
timestamp 1626908933
transform 1 0 6528 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_495
timestamp 1626908933
transform 1 0 6528 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_16
timestamp 1626908933
transform 1 0 6912 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_71
timestamp 1626908933
transform 1 0 6912 0 -1 11988
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1109
timestamp 1626908933
transform 1 0 7056 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_321
timestamp 1626908933
transform 1 0 7056 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1029
timestamp 1626908933
transform 1 0 7056 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_261
timestamp 1626908933
transform 1 0 7056 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1030
timestamp 1626908933
transform 1 0 7056 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_262
timestamp 1626908933
transform 1 0 7056 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_815
timestamp 1626908933
transform 1 0 7248 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_27
timestamp 1626908933
transform 1 0 7248 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1160
timestamp 1626908933
transform 1 0 7392 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_530
timestamp 1626908933
transform 1 0 7392 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_119
timestamp 1626908933
transform 1 0 7488 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_378
timestamp 1626908933
transform 1 0 7488 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_531
timestamp 1626908933
transform 1 0 7584 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1161
timestamp 1626908933
transform 1 0 7584 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_318
timestamp 1626908933
transform 1 0 7824 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1106
timestamp 1626908933
transform 1 0 7824 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_69
timestamp 1626908933
transform 1 0 7680 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_14
timestamp 1626908933
transform 1 0 7680 0 -1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_298
timestamp 1626908933
transform 1 0 8160 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_666
timestamp 1626908933
transform 1 0 8160 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_725
timestamp 1626908933
transform 1 0 8304 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1493
timestamp 1626908933
transform 1 0 8304 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_24
timestamp 1626908933
transform 1 0 8016 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_812
timestamp 1626908933
transform 1 0 8016 0 1 11655
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_366
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_96
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_366
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_96
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_366
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_96
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_103
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_391
timestamp 1626908933
transform 1 0 8600 0 1 11322
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1542
timestamp 1626908933
transform 1 0 8688 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_754
timestamp 1626908933
transform 1 0 8688 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_11
timestamp 1626908933
transform 1 0 8352 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_91
timestamp 1626908933
transform 1 0 8352 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_299
timestamp 1626908933
transform 1 0 9216 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_667
timestamp 1626908933
transform 1 0 9216 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_53
timestamp 1626908933
transform 1 0 8880 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_722
timestamp 1626908933
transform 1 0 8976 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_821
timestamp 1626908933
transform 1 0 8880 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1490
timestamp 1626908933
transform 1 0 8976 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_61
timestamp 1626908933
transform 1 0 9072 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_849
timestamp 1626908933
transform 1 0 9072 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_532
timestamp 1626908933
transform 1 0 9408 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1162
timestamp 1626908933
transform 1 0 9408 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_743
timestamp 1626908933
transform 1 0 9648 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1531
timestamp 1626908933
transform 1 0 9648 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_27
timestamp 1626908933
transform 1 0 9504 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_107
timestamp 1626908933
transform 1 0 9504 0 -1 11988
box -38 -49 902 715
use M1M2_PR  M1M2_PR_793
timestamp 1626908933
transform 1 0 9840 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_25
timestamp 1626908933
transform 1 0 9840 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_808
timestamp 1626908933
transform 1 0 10032 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_20
timestamp 1626908933
transform 1 0 10032 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1163
timestamp 1626908933
transform 1 0 10560 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_533
timestamp 1626908933
transform 1 0 10560 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_668
timestamp 1626908933
transform 1 0 10368 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_300
timestamp 1626908933
transform 1 0 10368 0 -1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_697
timestamp 1626908933
transform 1 0 10992 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1465
timestamp 1626908933
transform 1 0 10992 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_728
timestamp 1626908933
transform 1 0 10992 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1516
timestamp 1626908933
transform 1 0 10992 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_534
timestamp 1626908933
transform 1 0 11520 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1164
timestamp 1626908933
transform 1 0 11520 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_17
timestamp 1626908933
transform 1 0 11184 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_805
timestamp 1626908933
transform 1 0 11184 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_22
timestamp 1626908933
transform 1 0 10656 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_102
timestamp 1626908933
transform 1 0 10656 0 -1 11988
box -38 -49 902 715
use osc_core_VIA5  osc_core_VIA5_81
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_351
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_81
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_351
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_81
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_351
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_87
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_375
timestamp 1626908933
transform 1 0 12600 0 1 11322
box -200 -142 200 178
use M1M2_PR  M1M2_PR_20
timestamp 1626908933
transform 1 0 12336 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_788
timestamp 1626908933
transform 1 0 12336 0 1 11729
box -32 -32 32 32
use L1M1_PR  L1M1_PR_16
timestamp 1626908933
transform 1 0 12144 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_804
timestamp 1626908933
transform 1 0 12144 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_680
timestamp 1626908933
transform 1 0 11760 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1448
timestamp 1626908933
transform 1 0 11760 0 1 11655
box -32 -32 32 32
use L1M1_PR  L1M1_PR_713
timestamp 1626908933
transform 1 0 11760 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1501
timestamp 1626908933
transform 1 0 11760 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_18
timestamp 1626908933
transform 1 0 11616 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_98
timestamp 1626908933
transform 1 0 11616 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_118
timestamp 1626908933
transform 1 0 12480 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_377
timestamp 1626908933
transform 1 0 12480 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_396
timestamp 1626908933
transform 1 0 12672 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_965
timestamp 1626908933
transform 1 0 12672 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_154
timestamp 1626908933
transform 1 0 12576 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_784
timestamp 1626908933
transform 1 0 12576 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_673
timestamp 1626908933
transform 1 0 13104 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1441
timestamp 1626908933
transform 1 0 13104 0 1 11581
box -32 -32 32 32
use L1M1_PR  L1M1_PR_706
timestamp 1626908933
transform 1 0 13200 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1494
timestamp 1626908933
transform 1 0 13200 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_19
timestamp 1626908933
transform 1 0 13056 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_99
timestamp 1626908933
transform 1 0 13056 0 -1 11988
box -38 -49 902 715
use L1M1_PR  L1M1_PR_13
timestamp 1626908933
transform 1 0 13584 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_801
timestamp 1626908933
transform 1 0 13584 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_301
timestamp 1626908933
transform 1 0 13920 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_669
timestamp 1626908933
transform 1 0 13920 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_535
timestamp 1626908933
transform 1 0 14112 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1165
timestamp 1626908933
transform 1 0 14112 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_672
timestamp 1626908933
transform 1 0 14160 0 1 11137
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1440
timestamp 1626908933
transform 1 0 14160 0 1 11137
box -32 -32 32 32
use M1M2_PR  M1M2_PR_671
timestamp 1626908933
transform 1 0 14160 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1439
timestamp 1626908933
transform 1 0 14160 0 1 11581
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_16
timestamp 1626908933
transform 1 0 14208 0 -1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_96
timestamp 1626908933
transform 1 0 14208 0 -1 11988
box -38 -49 902 715
use L1M1_PR  L1M1_PR_6
timestamp 1626908933
transform 1 0 14736 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_702
timestamp 1626908933
transform 1 0 14352 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_794
timestamp 1626908933
transform 1 0 14736 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1490
timestamp 1626908933
transform 1 0 14352 0 1 11655
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_351
timestamp 1626908933
transform 1 0 15168 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_920
timestamp 1626908933
transform 1 0 15168 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_153
timestamp 1626908933
transform 1 0 15072 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_783
timestamp 1626908933
transform 1 0 15072 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_11
timestamp 1626908933
transform 1 0 14928 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_779
timestamp 1626908933
transform 1 0 14928 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_958
timestamp 1626908933
transform 1 0 15552 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_388
timestamp 1626908933
transform 1 0 15552 0 -1 11988
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_66
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_336
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_66
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_336
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_66
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_336
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_71
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_359
timestamp 1626908933
transform 1 0 16600 0 1 11322
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_326
timestamp 1626908933
transform 1 0 16320 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_895
timestamp 1626908933
transform 1 0 16320 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_362
timestamp 1626908933
transform 1 0 16704 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_932
timestamp 1626908933
transform 1 0 16704 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_376
timestamp 1626908933
transform 1 0 17472 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_117
timestamp 1626908933
transform 1 0 17472 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_470
timestamp 1626908933
transform 1 0 17568 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_102
timestamp 1626908933
transform 1 0 17568 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_870
timestamp 1626908933
transform 1 0 17760 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_301
timestamp 1626908933
transform 1 0 17760 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_909
timestamp 1626908933
transform 1 0 18144 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_339
timestamp 1626908933
transform 1 0 18144 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_853
timestamp 1626908933
transform 1 0 18912 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_284
timestamp 1626908933
transform 1 0 18912 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_782
timestamp 1626908933
transform 1 0 19296 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_152
timestamp 1626908933
transform 1 0 19296 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_887
timestamp 1626908933
transform 1 0 19392 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_317
timestamp 1626908933
transform 1 0 19392 0 -1 11988
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_321
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_51
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_321
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_51
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_321
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_51
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_55
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_343
timestamp 1626908933
transform 1 0 20600 0 1 11322
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_469
timestamp 1626908933
transform 1 0 20160 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_101
timestamp 1626908933
transform 1 0 20160 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_268
timestamp 1626908933
transform 1 0 20352 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_837
timestamp 1626908933
transform 1 0 20352 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_859
timestamp 1626908933
transform 1 0 20736 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_289
timestamp 1626908933
transform 1 0 20736 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_468
timestamp 1626908933
transform 1 0 21504 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_100
timestamp 1626908933
transform 1 0 21504 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_835
timestamp 1626908933
transform 1 0 21696 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_265
timestamp 1626908933
transform 1 0 21696 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_116
timestamp 1626908933
transform 1 0 22464 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_375
timestamp 1626908933
transform 1 0 22464 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_431
timestamp 1626908933
transform 1 0 22560 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1061
timestamp 1626908933
transform 1 0 22560 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_566
timestamp 1626908933
transform 1 0 22800 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1354
timestamp 1626908933
transform 1 0 22800 0 1 11729
box -29 -23 29 23
use M1M2_PR  M1M2_PR_464
timestamp 1626908933
transform 1 0 23280 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1232
timestamp 1626908933
transform 1 0 23280 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_496
timestamp 1626908933
transform 1 0 22896 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1264
timestamp 1626908933
transform 1 0 22896 0 1 11729
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_29
timestamp 1626908933
transform 1 0 22656 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_69
timestamp 1626908933
transform 1 0 22656 0 -1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1313
timestamp 1626908933
transform 1 0 23472 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_525
timestamp 1626908933
transform 1 0 23472 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_48
timestamp 1626908933
transform 1 0 23424 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_8
timestamp 1626908933
transform 1 0 23424 0 -1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_367
timestamp 1626908933
transform 1 0 23664 0 1 11063
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1135
timestamp 1626908933
transform 1 0 23664 0 1 11063
box -32 -32 32 32
use M1M2_PR  M1M2_PR_480
timestamp 1626908933
transform 1 0 24144 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1248
timestamp 1626908933
transform 1 0 24144 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_548
timestamp 1626908933
transform 1 0 24048 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1336
timestamp 1626908933
transform 1 0 24048 0 1 11211
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_36
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_306
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_36
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_306
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_36
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_306
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_327
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_39
timestamp 1626908933
transform 1 0 24600 0 1 11322
box -200 -142 200 178
use M1M2_PR  M1M2_PR_369
timestamp 1626908933
transform 1 0 24048 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1137
timestamp 1626908933
transform 1 0 24048 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1205
timestamp 1626908933
transform 1 0 25776 0 1 11507
box -32 -32 32 32
use M1M2_PR  M1M2_PR_437
timestamp 1626908933
transform 1 0 25776 0 1 11507
box -32 -32 32 32
use L1M1_PR  L1M1_PR_498
timestamp 1626908933
transform 1 0 26064 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1286
timestamp 1626908933
transform 1 0 26064 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_115
timestamp 1626908933
transform 1 0 26112 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_374
timestamp 1626908933
transform 1 0 26112 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_496
timestamp 1626908933
transform 1 0 25968 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1284
timestamp 1626908933
transform 1 0 25968 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_432
timestamp 1626908933
transform 1 0 26160 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1200
timestamp 1626908933
transform 1 0 26160 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_431
timestamp 1626908933
transform 1 0 26160 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1199
timestamp 1626908933
transform 1 0 26160 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_9
timestamp 1626908933
transform 1 0 25824 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_4
timestamp 1626908933
transform 1 0 25824 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_33
timestamp 1626908933
transform 1 0 26208 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_73
timestamp 1626908933
transform 1 0 26208 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_28
timestamp 1626908933
transform 1 0 24192 0 -1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_12
timestamp 1626908933
transform 1 0 24192 0 -1 11988
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_524
timestamp 1626908933
transform 1 0 27024 0 1 11211
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1292
timestamp 1626908933
transform 1 0 27024 0 1 11211
box -32 -32 32 32
use L1M1_PR  L1M1_PR_597
timestamp 1626908933
transform 1 0 27024 0 1 11211
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1385
timestamp 1626908933
transform 1 0 27024 0 1 11211
box -29 -23 29 23
use M1M2_PR  M1M2_PR_523
timestamp 1626908933
transform 1 0 27024 0 1 11581
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1291
timestamp 1626908933
transform 1 0 27024 0 1 11581
box -32 -32 32 32
use L1M1_PR  L1M1_PR_603
timestamp 1626908933
transform 1 0 26352 0 1 11729
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1391
timestamp 1626908933
transform 1 0 26352 0 1 11729
box -29 -23 29 23
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_13
timestamp 1626908933
transform 1 0 26976 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  sky130_fd_sc_hs__clkbuf_2_4
timestamp 1626908933
transform 1 0 26976 0 -1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1384
timestamp 1626908933
transform 1 0 27216 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_596
timestamp 1626908933
transform 1 0 27216 0 1 11581
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1276
timestamp 1626908933
transform 1 0 27504 0 1 11655
box -29 -23 29 23
use L1M1_PR  L1M1_PR_488
timestamp 1626908933
transform 1 0 27504 0 1 11655
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1186
timestamp 1626908933
transform 1 0 27504 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_418
timestamp 1626908933
transform 1 0 27504 0 1 11655
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_373
timestamp 1626908933
transform 1 0 27360 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_114
timestamp 1626908933
transform 1 0 27360 0 -1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1187
timestamp 1626908933
transform 1 0 27504 0 1 11433
box -32 -32 32 32
use M1M2_PR  M1M2_PR_419
timestamp 1626908933
transform 1 0 27504 0 1 11433
box -32 -32 32 32
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_7
timestamp 1626908933
transform 1 0 27456 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_2
timestamp 1626908933
transform 1 0 27456 0 -1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_151
timestamp 1626908933
transform 1 0 27744 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_781
timestamp 1626908933
transform 1 0 27744 0 -1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_489
timestamp 1626908933
transform 1 0 27696 0 1 11433
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1277
timestamp 1626908933
transform 1 0 27696 0 1 11433
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_161
timestamp 1626908933
transform 1 0 27840 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_731
timestamp 1626908933
transform 1 0 27840 0 -1 11988
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_311
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_23
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_291
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_21
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_291
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_21
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_291
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_21
timestamp 1626908933
transform 1 0 28600 0 1 11322
box -200 -49 200 49
use M1M2_PR  M1M2_PR_1149
timestamp 1626908933
transform 1 0 28656 0 1 11729
box -32 -32 32 32
use M1M2_PR  M1M2_PR_381
timestamp 1626908933
transform 1 0 28656 0 1 11729
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_467
timestamp 1626908933
transform 1 0 28608 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_99
timestamp 1626908933
transform 1 0 28608 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_150
timestamp 1626908933
transform 1 0 28800 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_780
timestamp 1626908933
transform 1 0 28800 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_707
timestamp 1626908933
transform 1 0 28896 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_137
timestamp 1626908933
transform 1 0 28896 0 -1 11988
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1147
timestamp 1626908933
transform 1 0 28848 0 1 11063
box -32 -32 32 32
use M1M2_PR  M1M2_PR_379
timestamp 1626908933
transform 1 0 28848 0 1 11063
box -32 -32 32 32
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_3
timestamp 1626908933
transform 1 0 29664 0 -1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_19
timestamp 1626908933
transform 1 0 29664 0 -1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_87
timestamp 1626908933
transform 1 0 31680 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_657
timestamp 1626908933
transform 1 0 31680 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_96
timestamp 1626908933
transform 1 0 31296 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_665
timestamp 1626908933
transform 1 0 31296 0 -1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_415
timestamp 1626908933
transform 1 0 29712 0 1 11655
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1183
timestamp 1626908933
transform 1 0 29712 0 1 11655
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_295
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_7
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_276
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_6
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_276
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_6
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_276
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_6
timestamp 1626908933
transform 1 0 32600 0 1 11322
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_372
timestamp 1626908933
transform 1 0 32448 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_113
timestamp 1626908933
transform 1 0 32448 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_63
timestamp 1626908933
transform 1 0 32544 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_632
timestamp 1626908933
transform 1 0 32544 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_627
timestamp 1626908933
transform 1 0 32928 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_57
timestamp 1626908933
transform 1 0 32928 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_779
timestamp 1626908933
transform 1 0 33696 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_149
timestamp 1626908933
transform 1 0 33696 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_599
timestamp 1626908933
transform 1 0 33792 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_30
timestamp 1626908933
transform 1 0 33792 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_597
timestamp 1626908933
transform 1 0 34176 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_27
timestamp 1626908933
transform 1 0 34176 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_6
timestamp 1626908933
transform 1 0 34944 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_576
timestamp 1626908933
transform 1 0 34944 0 -1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_685
timestamp 1626908933
transform 1 0 144 0 1 11803
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1473
timestamp 1626908933
transform 1 0 144 0 1 11803
box -29 -23 29 23
use M2M3_PR  M2M3_PR_50
timestamp 1626908933
transform 1 0 48 0 1 12359
box -33 -37 33 37
use M2M3_PR  M2M3_PR_109
timestamp 1626908933
transform 1 0 48 0 1 12359
box -33 -37 33 37
use M1M2_PR  M1M2_PR_652
timestamp 1626908933
transform 1 0 144 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1420
timestamp 1626908933
transform 1 0 144 0 1 12247
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_112
timestamp 1626908933
transform 1 0 288 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_371
timestamp 1626908933
transform 1 0 288 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_399
timestamp 1626908933
transform 1 0 336 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1167
timestamp 1626908933
transform 1 0 336 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_682
timestamp 1626908933
transform 1 0 432 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1470
timestamp 1626908933
transform 1 0 432 0 1 12247
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_6
timestamp 1626908933
transform 1 0 384 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_31
timestamp 1626908933
transform 1 0 384 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_269
timestamp 1626908933
transform 1 0 624 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1037
timestamp 1626908933
transform 1 0 624 0 1 12099
box -32 -32 32 32
use L1M1_PR  L1M1_PR_331
timestamp 1626908933
transform 1 0 624 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1119
timestamp 1626908933
transform 1 0 624 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_683
timestamp 1626908933
transform 1 0 912 0 1 11803
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1471
timestamp 1626908933
transform 1 0 912 0 1 11803
box -29 -23 29 23
use M1M2_PR  M1M2_PR_391
timestamp 1626908933
transform 1 0 912 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1159
timestamp 1626908933
transform 1 0 912 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_328
timestamp 1626908933
transform 1 0 720 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1096
timestamp 1626908933
transform 1 0 720 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_401
timestamp 1626908933
transform 1 0 720 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1189
timestamp 1626908933
transform 1 0 720 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_473
timestamp 1626908933
transform 1 0 528 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1261
timestamp 1626908933
transform 1 0 528 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_302
timestamp 1626908933
transform 1 0 768 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_670
timestamp 1626908933
transform 1 0 768 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_334
timestamp 1626908933
transform 1 0 1200 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_339
timestamp 1626908933
transform 1 0 1200 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1122
timestamp 1626908933
transform 1 0 1200 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1127
timestamp 1626908933
transform 1 0 1200 0 1 12099
box -29 -23 29 23
use M1M2_PR  M1M2_PR_333
timestamp 1626908933
transform 1 0 1104 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1101
timestamp 1626908933
transform 1 0 1104 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_336
timestamp 1626908933
transform 1 0 1296 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1104
timestamp 1626908933
transform 1 0 1296 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_413
timestamp 1626908933
transform 1 0 1296 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1201
timestamp 1626908933
transform 1 0 1296 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_462
timestamp 1626908933
transform 1 0 1104 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1250
timestamp 1626908933
transform 1 0 1104 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_303
timestamp 1626908933
transform 1 0 1344 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_671
timestamp 1626908933
transform 1 0 1344 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_8
timestamp 1626908933
transform 1 0 960 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_33
timestamp 1626908933
transform 1 0 960 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1042
timestamp 1626908933
transform 1 0 1488 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_274
timestamp 1626908933
transform 1 0 1488 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1092
timestamp 1626908933
transform 1 0 1680 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_324
timestamp 1626908933
transform 1 0 1680 0 1 11877
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1185
timestamp 1626908933
transform 1 0 1872 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_397
timestamp 1626908933
transform 1 0 1872 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1045
timestamp 1626908933
transform 1 0 1968 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_277
timestamp 1626908933
transform 1 0 1968 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1046
timestamp 1626908933
transform 1 0 1872 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_278
timestamp 1626908933
transform 1 0 1872 0 1 12099
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1134
timestamp 1626908933
transform 1 0 1776 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_346
timestamp 1626908933
transform 1 0 1776 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1052
timestamp 1626908933
transform 1 0 1776 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_284
timestamp 1626908933
transform 1 0 1776 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1476
timestamp 1626908933
transform 1 0 1872 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_688
timestamp 1626908933
transform 1 0 1872 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1424
timestamp 1626908933
transform 1 0 1872 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_656
timestamp 1626908933
transform 1 0 1872 0 1 12247
box -32 -32 32 32
use M2M3_PR  M2M3_PR_108
timestamp 1626908933
transform 1 0 1872 0 1 12359
box -33 -37 33 37
use M2M3_PR  M2M3_PR_49
timestamp 1626908933
transform 1 0 1872 0 1 12359
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1041
timestamp 1626908933
transform 1 0 1584 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_273
timestamp 1626908933
transform 1 0 1584 0 1 12469
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_18
timestamp 1626908933
transform 1 0 1824 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_43
timestamp 1626908933
transform 1 0 1824 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_3
timestamp 1626908933
transform -1 0 1824 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_8
timestamp 1626908933
transform -1 0 1824 0 1 11988
box -38 -49 326 715
use L1M1_PR  L1M1_PR_1475
timestamp 1626908933
transform 1 0 2064 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_687
timestamp 1626908933
transform 1 0 2064 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1423
timestamp 1626908933
transform 1 0 2064 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_655
timestamp 1626908933
transform 1 0 2064 0 1 11877
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1100
timestamp 1626908933
transform 1 0 2352 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_312
timestamp 1626908933
transform 1 0 2352 0 1 11877
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_531
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_261
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_531
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_261
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_531
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_261
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_566
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_278
timestamp 1626908933
transform 1 0 2600 0 1 11988
box -200 -142 200 178
use L1M1_PR  L1M1_PR_457
timestamp 1626908933
transform 1 0 1968 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1245
timestamp 1626908933
transform 1 0 1968 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_352
timestamp 1626908933
transform 1 0 2064 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1120
timestamp 1626908933
transform 1 0 2064 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_427
timestamp 1626908933
transform 1 0 2160 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1215
timestamp 1626908933
transform 1 0 2160 0 1 12247
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_78
timestamp 1626908933
transform 1 0 2496 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_23
timestamp 1626908933
transform 1 0 2496 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_536
timestamp 1626908933
transform 1 0 2400 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1166
timestamp 1626908933
transform 1 0 2400 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_304
timestamp 1626908933
transform 1 0 2208 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_672
timestamp 1626908933
transform 1 0 2208 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_901
timestamp 1626908933
transform 1 0 2832 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_113
timestamp 1626908933
transform 1 0 2832 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_865
timestamp 1626908933
transform 1 0 2832 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_97
timestamp 1626908933
transform 1 0 2832 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1121
timestamp 1626908933
transform 1 0 2640 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_333
timestamp 1626908933
transform 1 0 2640 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_4
timestamp 1626908933
transform 1 0 2976 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_59
timestamp 1626908933
transform 1 0 2976 0 1 11988
box -38 -49 518 715
use M1M2_PR  M1M2_PR_832
timestamp 1626908933
transform 1 0 3312 0 1 12173
box -32 -32 32 32
use M1M2_PR  M1M2_PR_64
timestamp 1626908933
transform 1 0 3312 0 1 12173
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1092
timestamp 1626908933
transform 1 0 3216 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_863
timestamp 1626908933
transform 1 0 3312 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_304
timestamp 1626908933
transform 1 0 3216 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_75
timestamp 1626908933
transform 1 0 3312 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1019
timestamp 1626908933
transform 1 0 3216 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_251
timestamp 1626908933
transform 1 0 3216 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1090
timestamp 1626908933
transform 1 0 3600 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_302
timestamp 1626908933
transform 1 0 3600 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1017
timestamp 1626908933
transform 1 0 3504 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_249
timestamp 1626908933
transform 1 0 3504 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_61
timestamp 1626908933
transform 1 0 3456 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_6
timestamp 1626908933
transform 1 0 3456 0 1 11988
box -38 -49 518 715
use L1M1_PR  L1M1_PR_860
timestamp 1626908933
transform 1 0 3792 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_72
timestamp 1626908933
transform 1 0 3792 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1167
timestamp 1626908933
transform 1 0 3936 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_537
timestamp 1626908933
transform 1 0 3936 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_26
timestamp 1626908933
transform 1 0 4032 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_81
timestamp 1626908933
transform 1 0 4032 0 1 11988
box -38 -49 518 715
use M1M2_PR  M1M2_PR_276
timestamp 1626908933
transform 1 0 4560 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1044
timestamp 1626908933
transform 1 0 4560 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_275
timestamp 1626908933
transform 1 0 4560 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1043
timestamp 1626908933
transform 1 0 4560 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_109
timestamp 1626908933
transform 1 0 4368 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_337
timestamp 1626908933
transform 1 0 4656 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_338
timestamp 1626908933
transform 1 0 4272 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_897
timestamp 1626908933
transform 1 0 4368 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1125
timestamp 1626908933
transform 1 0 4656 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1126
timestamp 1626908933
transform 1 0 4272 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_80
timestamp 1626908933
transform 1 0 4512 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_25
timestamp 1626908933
transform 1 0 4512 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_111
timestamp 1626908933
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_370
timestamp 1626908933
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_88
timestamp 1626908933
transform 1 0 4944 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_856
timestamp 1626908933
transform 1 0 4944 0 1 12395
box -32 -32 32 32
use L1M1_PR  L1M1_PR_102
timestamp 1626908933
transform 1 0 4848 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_890
timestamp 1626908933
transform 1 0 4848 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_335
timestamp 1626908933
transform 1 0 5232 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1123
timestamp 1626908933
transform 1 0 5232 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_82
timestamp 1626908933
transform 1 0 5088 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_27
timestamp 1626908933
transform 1 0 5088 0 1 11988
box -38 -49 518 715
use L1M1_PR  L1M1_PR_311
timestamp 1626908933
transform 1 0 5712 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1099
timestamp 1626908933
transform 1 0 5712 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_83
timestamp 1626908933
transform 1 0 5328 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_851
timestamp 1626908933
transform 1 0 5328 0 1 12395
box -32 -32 32 32
use L1M1_PR  L1M1_PR_97
timestamp 1626908933
transform 1 0 5424 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_885
timestamp 1626908933
transform 1 0 5424 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_255
timestamp 1626908933
transform 1 0 5616 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1023
timestamp 1626908933
transform 1 0 5616 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_508
timestamp 1626908933
transform 1 0 5568 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1077
timestamp 1626908933
transform 1 0 5568 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_35
timestamp 1626908933
transform 1 0 6192 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_803
timestamp 1626908933
transform 1 0 6192 0 1 11803
box -32 -32 32 32
use L1M1_PR  L1M1_PR_313
timestamp 1626908933
transform 1 0 6096 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1101
timestamp 1626908933
transform 1 0 6096 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_34
timestamp 1626908933
transform 1 0 6192 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_802
timestamp 1626908933
transform 1 0 6192 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_35
timestamp 1626908933
transform 1 0 6288 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_823
timestamp 1626908933
transform 1 0 6288 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_66
timestamp 1626908933
transform 1 0 5952 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_11
timestamp 1626908933
transform 1 0 5952 0 1 11988
box -38 -49 518 715
use osc_core_VIA5  osc_core_VIA5_246
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_516
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_246
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_516
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_246
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_516
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_262
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_550
timestamp 1626908933
transform 1 0 6600 0 1 11988
box -200 -142 200 178
use L1M1_PR  L1M1_PR_324
timestamp 1626908933
transform 1 0 6672 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1112
timestamp 1626908933
transform 1 0 6672 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_31
timestamp 1626908933
transform 1 0 6864 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_819
timestamp 1626908933
transform 1 0 6864 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_74
timestamp 1626908933
transform 1 0 6528 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_19
timestamp 1626908933
transform 1 0 6528 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_538
timestamp 1626908933
transform 1 0 6432 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1168
timestamp 1626908933
transform 1 0 6432 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_26
timestamp 1626908933
transform 1 0 7344 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_320
timestamp 1626908933
transform 1 0 7248 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_814
timestamp 1626908933
transform 1 0 7344 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1108
timestamp 1626908933
transform 1 0 7248 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_260
timestamp 1626908933
transform 1 0 7056 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1028
timestamp 1626908933
transform 1 0 7056 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_539
timestamp 1626908933
transform 1 0 7488 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1169
timestamp 1626908933
transform 1 0 7488 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_319
timestamp 1626908933
transform 1 0 7728 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1107
timestamp 1626908933
transform 1 0 7728 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_72
timestamp 1626908933
transform 1 0 7584 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_17
timestamp 1626908933
transform 1 0 7584 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_70
timestamp 1626908933
transform 1 0 7008 0 1 11988
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_15
timestamp 1626908933
transform 1 0 7008 0 1 11988
box -38 -49 518 715
use L1M1_PR  L1M1_PR_811
timestamp 1626908933
transform 1 0 8400 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_23
timestamp 1626908933
transform 1 0 8400 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_813
timestamp 1626908933
transform 1 0 7920 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_25
timestamp 1626908933
transform 1 0 7920 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_104
timestamp 1626908933
transform -1 0 9120 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_24
timestamp 1626908933
transform -1 0 9120 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_673
timestamp 1626908933
transform 1 0 8064 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_305
timestamp 1626908933
transform 1 0 8064 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1537
timestamp 1626908933
transform 1 0 9264 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_749
timestamp 1626908933
transform 1 0 9264 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1539
timestamp 1626908933
transform 1 0 8976 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_751
timestamp 1626908933
transform 1 0 8976 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1489
timestamp 1626908933
transform 1 0 8976 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_721
timestamp 1626908933
transform 1 0 8976 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_106
timestamp 1626908933
transform 1 0 9120 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_26
timestamp 1626908933
transform 1 0 9120 0 1 11988
box -38 -49 902 715
use L1M1_PR  L1M1_PR_810
timestamp 1626908933
transform 1 0 9840 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_22
timestamp 1626908933
transform 1 0 9840 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_792
timestamp 1626908933
transform 1 0 9840 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_24
timestamp 1626908933
transform 1 0 9840 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_778
timestamp 1626908933
transform 1 0 10080 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_148
timestamp 1626908933
transform 1 0 10080 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_369
timestamp 1626908933
transform 1 0 9984 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_110
timestamp 1626908933
transform 1 0 9984 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1015
timestamp 1626908933
transform 1 0 10176 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_446
timestamp 1626908933
transform 1 0 10176 0 1 11988
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_534
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_246
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_231
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_501
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_231
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_501
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_231
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_501
timestamp 1626908933
transform 1 0 10600 0 1 11988
box -200 -49 200 49
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_21
timestamp 1626908933
transform 1 0 10560 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_101
timestamp 1626908933
transform 1 0 10560 0 1 11988
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1517
timestamp 1626908933
transform 1 0 10800 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_806
timestamp 1626908933
transform 1 0 11088 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_729
timestamp 1626908933
transform 1 0 10800 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_18
timestamp 1626908933
transform 1 0 11088 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1464
timestamp 1626908933
transform 1 0 10992 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_696
timestamp 1626908933
transform 1 0 10992 0 1 12395
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_674
timestamp 1626908933
transform 1 0 11424 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_306
timestamp 1626908933
transform 1 0 11424 0 1 11988
box -38 -49 230 715
use M1M2_PR  M1M2_PR_679
timestamp 1626908933
transform 1 0 11760 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1447
timestamp 1626908933
transform 1 0 11760 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_712
timestamp 1626908933
transform 1 0 11760 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1500
timestamp 1626908933
transform 1 0 11760 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_74
timestamp 1626908933
transform 1 0 12144 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_842
timestamp 1626908933
transform 1 0 12144 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_84
timestamp 1626908933
transform 1 0 12144 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_872
timestamp 1626908933
transform 1 0 12144 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_34
timestamp 1626908933
transform 1 0 11616 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_114
timestamp 1626908933
transform 1 0 11616 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_995
timestamp 1626908933
transform 1 0 12960 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_425
timestamp 1626908933
transform 1 0 12960 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_777
timestamp 1626908933
transform 1 0 12864 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_147
timestamp 1626908933
transform 1 0 12864 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_974
timestamp 1626908933
transform 1 0 12480 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_405
timestamp 1626908933
transform 1 0 12480 0 1 11988
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1492
timestamp 1626908933
transform 1 0 14256 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_704
timestamp 1626908933
transform 1 0 14256 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1438
timestamp 1626908933
transform 1 0 14160 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_670
timestamp 1626908933
transform 1 0 14160 0 1 12247
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_97
timestamp 1626908933
transform 1 0 14112 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_17
timestamp 1626908933
transform 1 0 14112 0 1 11988
box -38 -49 902 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_942
timestamp 1626908933
transform 1 0 13728 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_373
timestamp 1626908933
transform 1 0 13728 0 1 11988
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_486
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_216
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_486
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_216
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_486
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_216
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_230
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_518
timestamp 1626908933
transform 1 0 14600 0 1 11988
box -200 -142 200 178
use L1M1_PR  L1M1_PR_798
timestamp 1626908933
transform 1 0 14640 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_10
timestamp 1626908933
transform 1 0 14640 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_783
timestamp 1626908933
transform 1 0 14640 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_15
timestamp 1626908933
transform 1 0 14640 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_109
timestamp 1626908933
transform 1 0 14976 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_368
timestamp 1626908933
transform 1 0 14976 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_350
timestamp 1626908933
transform 1 0 15168 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_919
timestamp 1626908933
transform 1 0 15168 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_146
timestamp 1626908933
transform 1 0 15072 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_776
timestamp 1626908933
transform 1 0 15072 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_957
timestamp 1626908933
transform 1 0 15552 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_387
timestamp 1626908933
transform 1 0 15552 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_931
timestamp 1626908933
transform 1 0 16704 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_361
timestamp 1626908933
transform 1 0 16704 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_894
timestamp 1626908933
transform 1 0 16320 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_325
timestamp 1626908933
transform 1 0 16320 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_367
timestamp 1626908933
transform 1 0 17472 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_108
timestamp 1626908933
transform 1 0 17472 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_466
timestamp 1626908933
transform 1 0 17568 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_98
timestamp 1626908933
transform 1 0 17568 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_869
timestamp 1626908933
transform 1 0 17760 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_300
timestamp 1626908933
transform 1 0 17760 0 1 11988
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_502
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_214
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_201
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_471
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_201
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_471
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_201
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_471
timestamp 1626908933
transform 1 0 18600 0 1 11988
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_338
timestamp 1626908933
transform 1 0 18144 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_908
timestamp 1626908933
transform 1 0 18144 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_775
timestamp 1626908933
transform 1 0 19104 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_145
timestamp 1626908933
transform 1 0 19104 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_465
timestamp 1626908933
transform 1 0 18912 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_97
timestamp 1626908933
transform 1 0 18912 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_886
timestamp 1626908933
transform 1 0 19200 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_316
timestamp 1626908933
transform 1 0 19200 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_870
timestamp 1626908933
transform 1 0 20064 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_300
timestamp 1626908933
transform 1 0 20064 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_366
timestamp 1626908933
transform 1 0 19968 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_107
timestamp 1626908933
transform 1 0 19968 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_464
timestamp 1626908933
transform 1 0 20832 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_96
timestamp 1626908933
transform 1 0 20832 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_821
timestamp 1626908933
transform 1 0 21024 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_252
timestamp 1626908933
transform 1 0 21024 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_844
timestamp 1626908933
transform 1 0 21408 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_274
timestamp 1626908933
transform 1 0 21408 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_95
timestamp 1626908933
transform 1 0 22176 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_463
timestamp 1626908933
transform 1 0 22176 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_540
timestamp 1626908933
transform 1 0 22368 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1170
timestamp 1626908933
transform 1 0 22368 0 1 11988
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_186
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_456
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_186
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_456
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_186
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_456
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_198
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_486
timestamp 1626908933
transform 1 0 22600 0 1 11988
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_106
timestamp 1626908933
transform 1 0 22464 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_365
timestamp 1626908933
transform 1 0 22464 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_532
timestamp 1626908933
transform 1 0 22608 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1320
timestamp 1626908933
transform 1 0 22608 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_463
timestamp 1626908933
transform 1 0 23280 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1231
timestamp 1626908933
transform 1 0 23280 0 1 12099
box -32 -32 32 32
use L1M1_PR  L1M1_PR_526
timestamp 1626908933
transform 1 0 23280 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1314
timestamp 1626908933
transform 1 0 23280 0 1 12099
box -29 -23 29 23
use M1M2_PR  M1M2_PR_492
timestamp 1626908933
transform 1 0 23184 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1260
timestamp 1626908933
transform 1 0 23184 0 1 11877
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_11
timestamp 1626908933
transform 1 0 22560 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_51
timestamp 1626908933
transform 1 0 22560 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1304
timestamp 1626908933
transform 1 0 23472 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_516
timestamp 1626908933
transform 1 0 23472 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_42
timestamp 1626908933
transform 1 0 23328 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_2
timestamp 1626908933
transform 1 0 23328 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1348
timestamp 1626908933
transform 1 0 23376 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_560
timestamp 1626908933
transform 1 0 23376 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_458
timestamp 1626908933
transform 1 0 23568 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1226
timestamp 1626908933
transform 1 0 23568 0 1 12321
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_105
timestamp 1626908933
transform 1 0 24096 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_364
timestamp 1626908933
transform 1 0 24096 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_520
timestamp 1626908933
transform 1 0 24144 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1308
timestamp 1626908933
transform 1 0 24144 0 1 11877
box -29 -23 29 23
use M1M2_PR  M1M2_PR_371
timestamp 1626908933
transform 1 0 24144 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_479
timestamp 1626908933
transform 1 0 24144 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1139
timestamp 1626908933
transform 1 0 24144 0 1 12395
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1247
timestamp 1626908933
transform 1 0 24144 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_500
timestamp 1626908933
transform 1 0 25584 0 1 11803
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1268
timestamp 1626908933
transform 1 0 25584 0 1 11803
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1283
timestamp 1626908933
transform 1 0 26064 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_495
timestamp 1626908933
transform 1 0 26064 0 1 12099
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1228
timestamp 1626908933
transform 1 0 25872 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1198
timestamp 1626908933
transform 1 0 26160 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_460
timestamp 1626908933
transform 1 0 25872 0 1 11877
box -32 -32 32 32
use M1M2_PR  M1M2_PR_430
timestamp 1626908933
transform 1 0 26160 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1204
timestamp 1626908933
transform 1 0 25776 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_436
timestamp 1626908933
transform 1 0 25776 0 1 12321
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1274
timestamp 1626908933
transform 1 0 25968 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_486
timestamp 1626908933
transform 1 0 25968 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1335
timestamp 1626908933
transform 1 0 26160 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_547
timestamp 1626908933
transform 1 0 26160 0 1 12247
box -29 -23 29 23
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_8
timestamp 1626908933
transform 1 0 25824 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_3
timestamp 1626908933
transform 1 0 25824 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_20
timestamp 1626908933
transform 1 0 26112 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_60
timestamp 1626908933
transform 1 0 26112 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_27
timestamp 1626908933
transform 1 0 24192 0 1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_11
timestamp 1626908933
transform 1 0 24192 0 1 11988
box -38 -49 1670 715
use osc_core_VIA4  osc_core_VIA4_182
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_470
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_171
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_441
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_171
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_441
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_171
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_441
timestamp 1626908933
transform 1 0 26600 0 1 11988
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_94
timestamp 1626908933
transform 1 0 26880 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_462
timestamp 1626908933
transform 1 0 26880 0 1 11988
box -38 -49 230 715
use L1M1_PR  L1M1_PR_571
timestamp 1626908933
transform 1 0 26928 0 1 11803
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1359
timestamp 1626908933
transform 1 0 26928 0 1 11803
box -29 -23 29 23
use L1M1_PR  L1M1_PR_602
timestamp 1626908933
transform 1 0 27120 0 1 11877
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1390
timestamp 1626908933
transform 1 0 27120 0 1 11877
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_170
timestamp 1626908933
transform 1 0 27072 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_739
timestamp 1626908933
transform 1 0 27072 0 1 11988
box -38 -49 422 715
use M1M2_PR  M1M2_PR_417
timestamp 1626908933
transform 1 0 27504 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1185
timestamp 1626908933
transform 1 0 27504 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_1
timestamp 1626908933
transform 1 0 27456 0 1 11988
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_6
timestamp 1626908933
transform 1 0 27456 0 1 11988
box -38 -49 326 715
use L1M1_PR  L1M1_PR_485
timestamp 1626908933
transform 1 0 27504 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1273
timestamp 1626908933
transform 1 0 27504 0 1 12321
box -29 -23 29 23
use M1M2_PR  M1M2_PR_466
timestamp 1626908933
transform 1 0 27408 0 1 12469
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1234
timestamp 1626908933
transform 1 0 27408 0 1 12469
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_144
timestamp 1626908933
transform 1 0 27744 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_774
timestamp 1626908933
transform 1 0 27744 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_487
timestamp 1626908933
transform 1 0 27696 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1275
timestamp 1626908933
transform 1 0 27696 0 1 12099
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_159
timestamp 1626908933
transform 1 0 27840 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_728
timestamp 1626908933
transform 1 0 27840 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_143
timestamp 1626908933
transform 1 0 28224 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_773
timestamp 1626908933
transform 1 0 28224 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_446
timestamp 1626908933
transform 1 0 28752 0 1 12099
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1234
timestamp 1626908933
transform 1 0 28752 0 1 12099
box -29 -23 29 23
use M1M2_PR  M1M2_PR_380
timestamp 1626908933
transform 1 0 28656 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1148
timestamp 1626908933
transform 1 0 28656 0 1 12247
box -32 -32 32 32
use L1M1_PR  L1M1_PR_447
timestamp 1626908933
transform 1 0 28656 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_484
timestamp 1626908933
transform 1 0 28464 0 1 12321
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1235
timestamp 1626908933
transform 1 0 28656 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1272
timestamp 1626908933
transform 1 0 28464 0 1 12321
box -29 -23 29 23
use sky130_fd_sc_hs__and4_2  sky130_fd_sc_hs__and4_2_0
timestamp 1626908933
transform -1 0 29088 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__and4_2  sky130_fd_sc_hs__and4_2_3
timestamp 1626908933
transform -1 0 29088 0 1 11988
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1237
timestamp 1626908933
transform 1 0 28848 0 1 12247
box -29 -23 29 23
use L1M1_PR  L1M1_PR_449
timestamp 1626908933
transform 1 0 28848 0 1 12247
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1146
timestamp 1626908933
transform 1 0 28848 0 1 12099
box -32 -32 32 32
use M1M2_PR  M1M2_PR_378
timestamp 1626908933
transform 1 0 28848 0 1 12099
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_131
timestamp 1626908933
transform 1 0 29184 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_700
timestamp 1626908933
transform 1 0 29184 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_142
timestamp 1626908933
transform 1 0 29088 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_772
timestamp 1626908933
transform 1 0 29088 0 1 11988
box -38 -49 134 715
use L1M1_PR  L1M1_PR_448
timestamp 1626908933
transform 1 0 29136 0 1 12395
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1236
timestamp 1626908933
transform 1 0 29136 0 1 12395
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_104
timestamp 1626908933
transform 1 0 29568 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_363
timestamp 1626908933
transform 1 0 29568 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_383
timestamp 1626908933
transform 1 0 29616 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_414
timestamp 1626908933
transform 1 0 29712 0 1 12321
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1151
timestamp 1626908933
transform 1 0 29616 0 1 12247
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1182
timestamp 1626908933
transform 1 0 29712 0 1 12321
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_454
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_166
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_156
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_426
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_156
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_426
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_156
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_426
timestamp 1626908933
transform 1 0 30600 0 1 11988
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_664
timestamp 1626908933
transform 1 0 31296 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_95
timestamp 1626908933
transform 1 0 31296 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_656
timestamp 1626908933
transform 1 0 31680 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_86
timestamp 1626908933
transform 1 0 31680 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_18
timestamp 1626908933
transform 1 0 29664 0 1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_2
timestamp 1626908933
transform 1 0 29664 0 1 11988
box -38 -49 1670 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_771
timestamp 1626908933
transform 1 0 32448 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_141
timestamp 1626908933
transform 1 0 32448 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_631
timestamp 1626908933
transform 1 0 32544 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_62
timestamp 1626908933
transform 1 0 32544 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_626
timestamp 1626908933
transform 1 0 32928 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_56
timestamp 1626908933
transform 1 0 32928 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_770
timestamp 1626908933
transform 1 0 33696 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_140
timestamp 1626908933
transform 1 0 33696 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_598
timestamp 1626908933
transform 1 0 33792 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_29
timestamp 1626908933
transform 1 0 33792 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_596
timestamp 1626908933
transform 1 0 34176 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_26
timestamp 1626908933
transform 1 0 34176 0 1 11988
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_411
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_141
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_411
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_141
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_411
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_141
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_150
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_438
timestamp 1626908933
transform 1 0 34600 0 1 11988
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_103
timestamp 1626908933
transform 1 0 34944 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_362
timestamp 1626908933
transform 1 0 34944 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_6
timestamp 1626908933
transform 1 0 35040 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_575
timestamp 1626908933
transform 1 0 35040 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_307
timestamp 1626908933
transform 1 0 35424 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_675
timestamp 1626908933
transform 1 0 35424 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_541
timestamp 1626908933
transform 1 0 35616 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1171
timestamp 1626908933
transform 1 0 35616 0 1 11988
box -38 -49 134 715
use M1M2_PR  M1M2_PR_654
timestamp 1626908933
transform 1 0 48 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1422
timestamp 1626908933
transform 1 0 48 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_653
timestamp 1626908933
transform 1 0 48 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1421
timestamp 1626908933
transform 1 0 48 0 1 13209
box -32 -32 32 32
use L1M1_PR  L1M1_PR_684
timestamp 1626908933
transform 1 0 144 0 1 13209
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1472
timestamp 1626908933
transform 1 0 144 0 1 13209
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_542
timestamp 1626908933
transform 1 0 288 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1172
timestamp 1626908933
transform 1 0 288 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_94
timestamp 1626908933
transform 1 0 288 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_353
timestamp 1626908933
transform 1 0 288 0 1 13320
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_395
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_125
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_395
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_125
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_395
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_125
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1136
timestamp 1626908933
transform 1 0 720 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_348
timestamp 1626908933
transform 1 0 720 0 1 12913
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_422
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_134
timestamp 1626908933
transform 1 0 600 0 1 12654
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1260
timestamp 1626908933
transform 1 0 528 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_472
timestamp 1626908933
transform 1 0 528 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1165
timestamp 1626908933
transform 1 0 528 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_397
timestamp 1626908933
transform 1 0 528 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1464
timestamp 1626908933
transform 1 0 432 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_676
timestamp 1626908933
transform 1 0 432 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1414
timestamp 1626908933
transform 1 0 336 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_646
timestamp 1626908933
transform 1 0 336 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1188
timestamp 1626908933
transform 1 0 720 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_400
timestamp 1626908933
transform 1 0 720 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1094
timestamp 1626908933
transform 1 0 816 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_326
timestamp 1626908933
transform 1 0 816 0 1 13061
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1176
timestamp 1626908933
transform 1 0 768 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_546
timestamp 1626908933
transform 1 0 768 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_29
timestamp 1626908933
transform 1 0 384 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_4
timestamp 1626908933
transform 1 0 384 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_38
timestamp 1626908933
transform 1 0 864 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_93
timestamp 1626908933
transform 1 0 864 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_28
timestamp 1626908933
transform 1 0 384 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_3
timestamp 1626908933
transform 1 0 384 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_33
timestamp 1626908933
transform 1 0 768 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_88
timestamp 1626908933
transform 1 0 768 0 -1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_686
timestamp 1626908933
transform 1 0 912 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1474
timestamp 1626908933
transform 1 0 912 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_195
timestamp 1626908933
transform 1 0 1104 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_347
timestamp 1626908933
transform 1 0 912 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_983
timestamp 1626908933
transform 1 0 1104 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1135
timestamp 1626908933
transform 1 0 912 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_286
timestamp 1626908933
transform 1 0 1296 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1054
timestamp 1626908933
transform 1 0 1296 0 1 12913
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_314
timestamp 1626908933
transform 1 0 1344 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_682
timestamp 1626908933
transform 1 0 1344 0 1 13320
box -38 -49 230 715
use L1M1_PR  L1M1_PR_350
timestamp 1626908933
transform 1 0 1392 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1138
timestamp 1626908933
transform 1 0 1392 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_90
timestamp 1626908933
transform 1 0 1248 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_35
timestamp 1626908933
transform 1 0 1248 0 -1 13320
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1091
timestamp 1626908933
transform 1 0 1680 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_323
timestamp 1626908933
transform 1 0 1680 0 1 12765
box -32 -32 32 32
use L1M1_PR  L1M1_PR_980
timestamp 1626908933
transform 1 0 1488 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_192
timestamp 1626908933
transform 1 0 1488 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_919
timestamp 1626908933
transform 1 0 1488 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_151
timestamp 1626908933
transform 1 0 1488 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_978
timestamp 1626908933
transform 1 0 1584 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_190
timestamp 1626908933
transform 1 0 1584 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_918
timestamp 1626908933
transform 1 0 1488 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_150
timestamp 1626908933
transform 1 0 1488 0 1 13061
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1137
timestamp 1626908933
transform 1 0 1872 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_349
timestamp 1626908933
transform 1 0 1872 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_46
timestamp 1626908933
transform 1 0 1536 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_21
timestamp 1626908933
transform 1 0 1536 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_13
timestamp 1626908933
transform 1 0 1920 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_4
timestamp 1626908933
transform 1 0 1920 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_34
timestamp 1626908933
transform 1 0 1728 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_89
timestamp 1626908933
transform 1 0 1728 0 -1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1115
timestamp 1626908933
transform 1 0 2256 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_327
timestamp 1626908933
transform 1 0 2256 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1040
timestamp 1626908933
transform 1 0 2064 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_272
timestamp 1626908933
transform 1 0 2064 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_187
timestamp 1626908933
transform 1 0 2064 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_975
timestamp 1626908933
transform 1 0 2064 0 1 12987
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_260
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_530
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_260
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_530
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_260
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_530
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_565
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_277
timestamp 1626908933
transform 1 0 2600 0 1 13320
box -200 -142 200 178
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_7
timestamp 1626908933
transform 1 0 2304 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_2
timestamp 1626908933
transform 1 0 2304 0 1 13320
box -38 -49 326 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_676
timestamp 1626908933
transform 1 0 2208 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_308
timestamp 1626908933
transform 1 0 2208 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1173
timestamp 1626908933
transform 1 0 2400 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_543
timestamp 1626908933
transform 1 0 2400 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_361
timestamp 1626908933
transform 1 0 2496 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_102
timestamp 1626908933
transform 1 0 2496 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_139
timestamp 1626908933
transform 1 0 2592 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_769
timestamp 1626908933
transform 1 0 2592 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_540
timestamp 1626908933
transform 1 0 2688 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1109
timestamp 1626908933
transform 1 0 2688 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_79
timestamp 1626908933
transform 1 0 2592 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_24
timestamp 1626908933
transform 1 0 2592 0 1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_396
timestamp 1626908933
transform 1 0 3120 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1184
timestamp 1626908933
transform 1 0 3120 0 1 12765
box -29 -23 29 23
use M3M4_PR  M3M4_PR_39
timestamp 1626908933
transform 1 0 3552 0 1 12969
box -38 -33 38 33
use M3M4_PR  M3M4_PR_18
timestamp 1626908933
transform 1 0 3552 0 1 12969
box -38 -33 38 33
use M2M3_PR  M2M3_PR_78
timestamp 1626908933
transform 1 0 3600 0 1 12969
box -33 -37 33 37
use M2M3_PR  M2M3_PR_19
timestamp 1626908933
transform 1 0 3600 0 1 12969
box -33 -37 33 37
use L1M1_PR  L1M1_PR_973
timestamp 1626908933
transform 1 0 3600 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_185
timestamp 1626908933
transform 1 0 3600 0 1 12913
box -29 -23 29 23
use M1M2_PR  M1M2_PR_916
timestamp 1626908933
transform 1 0 3600 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_148
timestamp 1626908933
transform 1 0 3600 0 1 12913
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1183
timestamp 1626908933
transform 1 0 3504 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_395
timestamp 1626908933
transform 1 0 3504 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1090
timestamp 1626908933
transform 1 0 3504 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_322
timestamp 1626908933
transform 1 0 3504 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_28
timestamp 1626908933
transform 1 0 3072 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_3
timestamp 1626908933
transform 1 0 3072 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_29
timestamp 1626908933
transform 1 0 3072 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_4
timestamp 1626908933
transform 1 0 3072 0 -1 13320
box -38 -49 1670 715
use osc_core_VIA4  osc_core_VIA4_118
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_406
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_380
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_110
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_380
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_110
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_380
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_110
timestamp 1626908933
transform 1 0 4600 0 1 12654
box -200 -49 200 49
use L1M1_PR  L1M1_PR_894
timestamp 1626908933
transform 1 0 4560 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_106
timestamp 1626908933
transform 1 0 4560 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_855
timestamp 1626908933
transform 1 0 4944 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_87
timestamp 1626908933
transform 1 0 4944 0 1 13061
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1177
timestamp 1626908933
transform 1 0 4896 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_547
timestamp 1626908933
transform 1 0 4896 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_352
timestamp 1626908933
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_93
timestamp 1626908933
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1174
timestamp 1626908933
transform 1 0 4896 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_544
timestamp 1626908933
transform 1 0 4896 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_683
timestamp 1626908933
transform 1 0 4704 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_315
timestamp 1626908933
transform 1 0 4704 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_677
timestamp 1626908933
transform 1 0 4704 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_309
timestamp 1626908933
transform 1 0 4704 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_86
timestamp 1626908933
transform 1 0 4992 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_31
timestamp 1626908933
transform 1 0 4992 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_87
timestamp 1626908933
transform 1 0 5088 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_32
timestamp 1626908933
transform 1 0 5088 0 1 13320
box -38 -49 518 715
use L1M1_PR  L1M1_PR_887
timestamp 1626908933
transform 1 0 5328 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_99
timestamp 1626908933
transform 1 0 5328 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1131
timestamp 1626908933
transform 1 0 5136 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_343
timestamp 1626908933
transform 1 0 5136 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1050
timestamp 1626908933
transform 1 0 5136 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_282
timestamp 1626908933
transform 1 0 5136 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_684
timestamp 1626908933
transform 1 0 5568 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_316
timestamp 1626908933
transform 1 0 5568 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1076
timestamp 1626908933
transform 1 0 5472 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_507
timestamp 1626908933
transform 1 0 5472 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1178
timestamp 1626908933
transform 1 0 5760 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_548
timestamp 1626908933
transform 1 0 5760 0 1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1114
timestamp 1626908933
transform 1 0 6000 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_326
timestamp 1626908933
transform 1 0 6000 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1034
timestamp 1626908933
transform 1 0 6000 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_266
timestamp 1626908933
transform 1 0 6000 0 1 12543
box -32 -32 32 32
use M2M3_PR  M2M3_PR_82
timestamp 1626908933
transform 1 0 6000 0 1 12969
box -33 -37 33 37
use M2M3_PR  M2M3_PR_23
timestamp 1626908933
transform 1 0 6000 0 1 12969
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1033
timestamp 1626908933
transform 1 0 6000 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_265
timestamp 1626908933
transform 1 0 6000 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_73
timestamp 1626908933
transform 1 0 5856 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_18
timestamp 1626908933
transform 1 0 5856 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_75
timestamp 1626908933
transform 1 0 5856 0 1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_20
timestamp 1626908933
transform 1 0 5856 0 1 13320
box -38 -49 518 715
use M1M2_PR  M1M2_PR_33
timestamp 1626908933
transform 1 0 6192 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_801
timestamp 1626908933
transform 1 0 6192 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_38
timestamp 1626908933
transform 1 0 6192 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_826
timestamp 1626908933
transform 1 0 6192 0 1 12987
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_245
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_515
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_245
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_515
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_245
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_515
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_549
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_261
timestamp 1626908933
transform 1 0 6600 0 1 13320
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1179
timestamp 1626908933
transform 1 0 6528 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_549
timestamp 1626908933
transform 1 0 6528 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_685
timestamp 1626908933
transform 1 0 6336 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_317
timestamp 1626908933
transform 1 0 6336 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_678
timestamp 1626908933
transform 1 0 6336 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_310
timestamp 1626908933
transform 1 0 6336 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_263
timestamp 1626908933
transform 1 0 6672 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1031
timestamp 1626908933
transform 1 0 6672 0 1 12987
box -32 -32 32 32
use M2M3_PR  M2M3_PR_22
timestamp 1626908933
transform 1 0 6672 0 1 12969
box -33 -37 33 37
use M2M3_PR  M2M3_PR_81
timestamp 1626908933
transform 1 0 6672 0 1 12969
box -33 -37 33 37
use L1M1_PR  L1M1_PR_30
timestamp 1626908933
transform 1 0 6864 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_323
timestamp 1626908933
transform 1 0 6672 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_818
timestamp 1626908933
transform 1 0 6864 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1111
timestamp 1626908933
transform 1 0 6672 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_76
timestamp 1626908933
transform 1 0 6528 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_21
timestamp 1626908933
transform 1 0 6528 0 -1 13320
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_30
timestamp 1626908933
transform 1 0 6624 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_110
timestamp 1626908933
transform 1 0 6624 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_491
timestamp 1626908933
transform 1 0 7104 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1060
timestamp 1626908933
transform 1 0 7104 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_138
timestamp 1626908933
transform 1 0 7008 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_768
timestamp 1626908933
transform 1 0 7008 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_101
timestamp 1626908933
transform 1 0 7488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_360
timestamp 1626908933
transform 1 0 7488 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_550
timestamp 1626908933
transform 1 0 7488 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1180
timestamp 1626908933
transform 1 0 7488 0 1 13320
box -38 -49 134 715
use M3M4_PR  M3M4_PR_31
timestamp 1626908933
transform 1 0 8112 0 1 12969
box -38 -33 38 33
use M3M4_PR  M3M4_PR_10
timestamp 1626908933
transform 1 0 8112 0 1 12969
box -38 -33 38 33
use M2M3_PR  M2M3_PR_70
timestamp 1626908933
transform 1 0 8112 0 1 12969
box -33 -37 33 37
use M2M3_PR  M2M3_PR_11
timestamp 1626908933
transform 1 0 8112 0 1 12969
box -33 -37 33 37
use L1M1_PR  L1M1_PR_920
timestamp 1626908933
transform 1 0 8112 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_132
timestamp 1626908933
transform 1 0 8112 0 1 12913
box -29 -23 29 23
use M1M2_PR  M1M2_PR_881
timestamp 1626908933
transform 1 0 8112 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_113
timestamp 1626908933
transform 1 0 8112 0 1 12913
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1176
timestamp 1626908933
transform 1 0 8304 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_388
timestamp 1626908933
transform 1 0 8304 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1085
timestamp 1626908933
transform 1 0 8304 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_317
timestamp 1626908933
transform 1 0 8304 0 1 12987
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_365
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_95
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_365
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_95
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_365
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_95
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_390
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_102
timestamp 1626908933
transform 1 0 8600 0 1 12654
box -200 -142 200 178
use L1M1_PR  L1M1_PR_955
timestamp 1626908933
transform 1 0 8976 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_167
timestamp 1626908933
transform 1 0 8976 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_901
timestamp 1626908933
transform 1 0 8976 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_133
timestamp 1626908933
transform 1 0 8976 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_455
timestamp 1626908933
transform 1 0 9216 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_87
timestamp 1626908933
transform 1 0 9216 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1175
timestamp 1626908933
transform 1 0 9216 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_545
timestamp 1626908933
transform 1 0 9216 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1488
timestamp 1626908933
transform 1 0 9072 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_720
timestamp 1626908933
transform 1 0 9072 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1533
timestamp 1626908933
transform 1 0 9456 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_745
timestamp 1626908933
transform 1 0 9456 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_760
timestamp 1626908933
transform 1 0 9408 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_130
timestamp 1626908933
transform 1 0 9408 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1033
timestamp 1626908933
transform 1 0 9504 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_464
timestamp 1626908933
transform 1 0 9504 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_25
timestamp 1626908933
transform 1 0 9312 0 -1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_105
timestamp 1626908933
transform 1 0 9312 0 -1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_48
timestamp 1626908933
transform 1 0 7584 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_23
timestamp 1626908933
transform 1 0 7584 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_49
timestamp 1626908933
transform 1 0 7584 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_24
timestamp 1626908933
transform 1 0 7584 0 -1 13320
box -38 -49 1670 715
use L1M1_PR  L1M1_PR_809
timestamp 1626908933
transform 1 0 9840 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_21
timestamp 1626908933
transform 1 0 9840 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_759
timestamp 1626908933
transform 1 0 9888 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_129
timestamp 1626908933
transform 1 0 9888 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_791
timestamp 1626908933
transform 1 0 9840 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_23
timestamp 1626908933
transform 1 0 9840 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_351
timestamp 1626908933
transform 1 0 9984 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_92
timestamp 1626908933
transform 1 0 9984 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_686
timestamp 1626908933
transform 1 0 10080 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_318
timestamp 1626908933
transform 1 0 10080 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_679
timestamp 1626908933
transform 1 0 10176 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_311
timestamp 1626908933
transform 1 0 10176 0 -1 13320
box -38 -49 230 715
use L1M1_PR  L1M1_PR_807
timestamp 1626908933
transform 1 0 10512 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_19
timestamp 1626908933
transform 1 0 10512 0 1 12987
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_245
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_533
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_500
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_230
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_500
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_230
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_500
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_230
timestamp 1626908933
transform 1 0 10600 0 1 13320
box -200 -49 200 49
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_23
timestamp 1626908933
transform -1 0 11232 0 -1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_103
timestamp 1626908933
transform -1 0 11232 0 -1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_48
timestamp 1626908933
transform 1 0 10272 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_128
timestamp 1626908933
transform 1 0 10272 0 1 13320
box -38 -49 902 715
use M1M2_PR  M1M2_PR_695
timestamp 1626908933
transform 1 0 10992 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1463
timestamp 1626908933
transform 1 0 10992 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_727
timestamp 1626908933
transform 1 0 10992 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1515
timestamp 1626908933
transform 1 0 10992 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_312
timestamp 1626908933
transform 1 0 11232 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_680
timestamp 1626908933
transform 1 0 11232 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_423
timestamp 1626908933
transform 1 0 11232 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_992
timestamp 1626908933
transform 1 0 11232 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_128
timestamp 1626908933
transform 1 0 11136 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_758
timestamp 1626908933
transform 1 0 11136 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_35
timestamp 1626908933
transform 1 0 11424 0 -1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_115
timestamp 1626908933
transform 1 0 11424 0 -1 13320
box -38 -49 902 715
use M1M2_PR  M1M2_PR_678
timestamp 1626908933
transform 1 0 11760 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1446
timestamp 1626908933
transform 1 0 11760 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_711
timestamp 1626908933
transform 1 0 11760 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1499
timestamp 1626908933
transform 1 0 11760 0 1 12987
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_80
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_350
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_80
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_350
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_80
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_350
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -49 200 49
use M2M3_PR  M2M3_PR_5
timestamp 1626908933
transform 1 0 12144 0 1 12847
box -33 -37 33 37
use M2M3_PR  M2M3_PR_64
timestamp 1626908933
transform 1 0 12144 0 1 12847
box -33 -37 33 37
use osc_core_VIA4  osc_core_VIA4_86
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_374
timestamp 1626908933
transform 1 0 12600 0 1 12654
box -200 -142 200 178
use L1M1_PR  L1M1_PR_871
timestamp 1626908933
transform 1 0 12144 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_83
timestamp 1626908933
transform 1 0 12144 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_841
timestamp 1626908933
transform 1 0 12144 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_73
timestamp 1626908933
transform 1 0 12144 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_681
timestamp 1626908933
transform 1 0 12288 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_313
timestamp 1626908933
transform 1 0 12288 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_32
timestamp 1626908933
transform 1 0 11616 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_112
timestamp 1626908933
transform 1 0 11616 0 1 13320
box -38 -49 902 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_359
timestamp 1626908933
transform 1 0 12480 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_100
timestamp 1626908933
transform 1 0 12480 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_973
timestamp 1626908933
transform 1 0 12480 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_404
timestamp 1626908933
transform 1 0 12480 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_687
timestamp 1626908933
transform 1 0 12864 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_319
timestamp 1626908933
transform 1 0 12864 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_461
timestamp 1626908933
transform 1 0 12576 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_93
timestamp 1626908933
transform 1 0 12576 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_964
timestamp 1626908933
transform 1 0 12768 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_395
timestamp 1626908933
transform 1 0 12768 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_551
timestamp 1626908933
transform 1 0 13056 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1181
timestamp 1626908933
transform 1 0 13056 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_311
timestamp 1626908933
transform 1 0 13680 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1079
timestamp 1626908933
transform 1 0 13680 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_383
timestamp 1626908933
transform 1 0 13680 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1171
timestamp 1626908933
transform 1 0 13680 0 1 12987
box -29 -23 29 23
use M3M4_PR  M3M4_PR_27
timestamp 1626908933
transform 1 0 14112 0 1 12847
box -38 -33 38 33
use M3M4_PR  M3M4_PR_6
timestamp 1626908933
transform 1 0 14112 0 1 12847
box -38 -33 38 33
use osc_core_VIA3  osc_core_VIA3_9
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_4
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_9
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_4
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -28 96 28
use osc_core_VIA1  osc_core_VIA1_9
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_4
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_9
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_4
timestamp 1626908933
transform 1 0 14116 0 1 13138
box -97 -33 96 33
use osc_core_VIA4  osc_core_VIA4_229
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_517
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_485
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_215
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_485
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_215
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_485
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_215
timestamp 1626908933
transform 1 0 14600 0 1 13320
box -200 -49 200 49
use L1M1_PR  L1M1_PR_797
timestamp 1626908933
transform 1 0 14640 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_9
timestamp 1626908933
transform 1 0 14640 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_688
timestamp 1626908933
transform 1 0 14784 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_320
timestamp 1626908933
transform 1 0 14784 0 1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_782
timestamp 1626908933
transform 1 0 14640 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_14
timestamp 1626908933
transform 1 0 14640 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_460
timestamp 1626908933
transform 1 0 14784 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_92
timestamp 1626908933
transform 1 0 14784 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_757
timestamp 1626908933
transform 1 0 15072 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_127
timestamp 1626908933
transform 1 0 15072 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_350
timestamp 1626908933
transform 1 0 14976 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_91
timestamp 1626908933
transform 1 0 14976 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_918
timestamp 1626908933
transform 1 0 15168 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_349
timestamp 1626908933
transform 1 0 15168 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_408
timestamp 1626908933
transform 1 0 14976 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_978
timestamp 1626908933
transform 1 0 14976 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_33
timestamp 1626908933
transform 1 0 13152 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_8
timestamp 1626908933
transform 1 0 13152 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_34
timestamp 1626908933
transform 1 0 13152 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_9
timestamp 1626908933
transform 1 0 13152 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_344
timestamp 1626908933
transform 1 0 15840 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_913
timestamp 1626908933
transform 1 0 15840 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_137
timestamp 1626908933
transform 1 0 15744 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_767
timestamp 1626908933
transform 1 0 15744 0 -1 13320
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_358
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_70
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_335
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_65
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_335
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_65
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_335
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_65
timestamp 1626908933
transform 1 0 16600 0 1 12654
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_893
timestamp 1626908933
transform 1 0 16320 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_324
timestamp 1626908933
transform 1 0 16320 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_379
timestamp 1626908933
transform 1 0 16224 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_949
timestamp 1626908933
transform 1 0 16224 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_386
timestamp 1626908933
transform 1 0 15552 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_956
timestamp 1626908933
transform 1 0 15552 0 1 13320
box -38 -49 806 715
use M1M2_PR  M1M2_PR_815
timestamp 1626908933
transform 1 0 18000 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_47
timestamp 1626908933
transform 1 0 18000 0 1 13209
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_930
timestamp 1626908933
transform 1 0 16704 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_360
timestamp 1626908933
transform 1 0 16704 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_889
timestamp 1626908933
transform 1 0 16992 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_320
timestamp 1626908933
transform 1 0 16992 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_358
timestamp 1626908933
transform 1 0 17376 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_99
timestamp 1626908933
transform 1 0 17376 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_43
timestamp 1626908933
transform 1 0 17472 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_18
timestamp 1626908933
transform 1 0 17472 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_44
timestamp 1626908933
transform 1 0 17472 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_19
timestamp 1626908933
transform 1 0 17472 0 -1 13320
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_548
timestamp 1626908933
transform 1 0 18288 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1316
timestamp 1626908933
transform 1 0 18288 0 1 12987
box -32 -32 32 32
use L1M1_PR  L1M1_PR_48
timestamp 1626908933
transform 1 0 18384 0 1 13135
box -29 -23 29 23
use L1M1_PR  L1M1_PR_623
timestamp 1626908933
transform 1 0 18288 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_836
timestamp 1626908933
transform 1 0 18384 0 1 13135
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1411
timestamp 1626908933
transform 1 0 18288 0 1 12987
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_213
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_501
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_200
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_470
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_200
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_470
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_200
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_470
timestamp 1626908933
transform 1 0 18600 0 1 13320
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_91
timestamp 1626908933
transform 1 0 19104 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_459
timestamp 1626908933
transform 1 0 19104 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_100
timestamp 1626908933
transform 1 0 19152 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_868
timestamp 1626908933
transform 1 0 19152 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_126
timestamp 1626908933
transform 1 0 19104 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_756
timestamp 1626908933
transform 1 0 19104 0 1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_118
timestamp 1626908933
transform 1 0 18960 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_906
timestamp 1626908933
transform 1 0 18960 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_136
timestamp 1626908933
transform 1 0 19296 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_766
timestamp 1626908933
transform 1 0 19296 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_315
timestamp 1626908933
transform 1 0 19392 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_885
timestamp 1626908933
transform 1 0 19392 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_314
timestamp 1626908933
transform 1 0 19200 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_884
timestamp 1626908933
transform 1 0 19200 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_90
timestamp 1626908933
transform 1 0 19968 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_349
timestamp 1626908933
transform 1 0 19968 0 1 13320
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_342
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_54
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_320
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_50
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_320
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_50
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_320
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_50
timestamp 1626908933
transform 1 0 20600 0 1 12654
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_765
timestamp 1626908933
transform 1 0 20160 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_135
timestamp 1626908933
transform 1 0 20160 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_267
timestamp 1626908933
transform 1 0 20256 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_836
timestamp 1626908933
transform 1 0 20256 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_299
timestamp 1626908933
transform 1 0 20064 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_869
timestamp 1626908933
transform 1 0 20064 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_858
timestamp 1626908933
transform 1 0 20640 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_288
timestamp 1626908933
transform 1 0 20640 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_251
timestamp 1626908933
transform 1 0 21120 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_820
timestamp 1626908933
transform 1 0 21120 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_86
timestamp 1626908933
transform 1 0 20832 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_454
timestamp 1626908933
transform 1 0 20832 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_125
timestamp 1626908933
transform 1 0 21024 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_755
timestamp 1626908933
transform 1 0 21024 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_98
timestamp 1626908933
transform 1 0 21408 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_357
timestamp 1626908933
transform 1 0 21408 0 -1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_554
timestamp 1626908933
transform 1 0 21936 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1322
timestamp 1626908933
transform 1 0 21936 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_597
timestamp 1626908933
transform 1 0 21744 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1365
timestamp 1626908933
transform 1 0 21744 0 1 13209
box -32 -32 32 32
use L1M1_PR  L1M1_PR_630
timestamp 1626908933
transform 1 0 21936 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1418
timestamp 1626908933
transform 1 0 21936 0 1 12987
box -29 -23 29 23
use M3M4_PR  M3M4_PR_22
timestamp 1626908933
transform 1 0 22224 0 1 13091
box -38 -33 38 33
use M3M4_PR  M3M4_PR_1
timestamp 1626908933
transform 1 0 22224 0 1 13091
box -38 -33 38 33
use M2M3_PR  M2M3_PR_59
timestamp 1626908933
transform 1 0 22416 0 1 13091
box -33 -37 33 37
use M2M3_PR  M2M3_PR_0
timestamp 1626908933
transform 1 0 22416 0 1 13091
box -33 -37 33 37
use L1M1_PR  L1M1_PR_790
timestamp 1626908933
transform 1 0 22416 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2
timestamp 1626908933
transform 1 0 22416 0 1 13061
box -29 -23 29 23
use M1M2_PR  M1M2_PR_768
timestamp 1626908933
transform 1 0 22416 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_0
timestamp 1626908933
transform 1 0 22416 0 1 13061
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_455
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_185
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_455
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_185
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_455
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_185
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_485
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_197
timestamp 1626908933
transform 1 0 22600 0 1 13320
box -200 -142 200 178
use L1M1_PR  L1M1_PR_831
timestamp 1626908933
transform 1 0 22992 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_43
timestamp 1626908933
transform 1 0 22992 0 1 12987
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_689
timestamp 1626908933
transform 1 0 23136 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_321
timestamp 1626908933
transform 1 0 23136 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_458
timestamp 1626908933
transform 1 0 23136 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_90
timestamp 1626908933
transform 1 0 23136 0 -1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_808
timestamp 1626908933
transform 1 0 22992 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_40
timestamp 1626908933
transform 1 0 22992 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_764
timestamp 1626908933
transform 1 0 23328 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_134
timestamp 1626908933
transform 1 0 23328 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_784
timestamp 1626908933
transform 1 0 23424 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_215
timestamp 1626908933
transform 1 0 23424 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__and4_2  sky130_fd_sc_hs__and4_2_2
timestamp 1626908933
transform -1 0 24096 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__and4_2  sky130_fd_sc_hs__and4_2_5
timestamp 1626908933
transform -1 0 24096 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_38
timestamp 1626908933
transform 1 0 21504 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_13
timestamp 1626908933
transform 1 0 21504 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_39
timestamp 1626908933
transform 1 0 21504 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_14
timestamp 1626908933
transform 1 0 21504 0 -1 13320
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_457
timestamp 1626908933
transform 1 0 23568 0 1 12839
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1225
timestamp 1626908933
transform 1 0 23568 0 1 12839
box -32 -32 32 32
use sky130_fd_sc_hs__clkbuf_1  sky130_fd_sc_hs__clkbuf_1_0
timestamp 1626908933
transform 1 0 23808 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  sky130_fd_sc_hs__clkbuf_1_1
timestamp 1626908933
transform 1 0 23808 0 -1 13320
box -38 -49 422 715
use L1M1_PR  L1M1_PR_508
timestamp 1626908933
transform 1 0 23952 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1296
timestamp 1626908933
transform 1 0 23952 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1295
timestamp 1626908933
transform 1 0 24048 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_507
timestamp 1626908933
transform 1 0 24048 0 1 12543
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1218
timestamp 1626908933
transform 1 0 24240 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_450
timestamp 1626908933
transform 1 0 24240 0 1 12543
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_305
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_35
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_305
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_35
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_305
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_35
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -49 200 49
use L1M1_PR  L1M1_PR_619
timestamp 1626908933
transform 1 0 24144 0 1 12913
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1407
timestamp 1626908933
transform 1 0 24144 0 1 12913
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_38
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_326
timestamp 1626908933
transform 1 0 24600 0 1 12654
box -200 -142 200 178
use M1M2_PR  M1M2_PR_1217
timestamp 1626908933
transform 1 0 24240 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_449
timestamp 1626908933
transform 1 0 24240 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_348
timestamp 1626908933
transform 1 0 24096 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_89
timestamp 1626908933
transform 1 0 24096 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_595
timestamp 1626908933
transform 1 0 25008 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1363
timestamp 1626908933
transform 1 0 25008 0 1 13209
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1238
timestamp 1626908933
transform 1 0 25776 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1211
timestamp 1626908933
transform 1 0 25680 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_470
timestamp 1626908933
transform 1 0 25776 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_443
timestamp 1626908933
transform 1 0 25680 0 1 13061
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1227
timestamp 1626908933
transform 1 0 25872 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_459
timestamp 1626908933
transform 1 0 25872 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_356
timestamp 1626908933
transform 1 0 25824 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_97
timestamp 1626908933
transform 1 0 25824 0 -1 13320
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1307
timestamp 1626908933
transform 1 0 25968 0 1 12987
box -29 -23 29 23
use L1M1_PR  L1M1_PR_519
timestamp 1626908933
transform 1 0 25968 0 1 12987
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1273
timestamp 1626908933
transform 1 0 26256 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_505
timestamp 1626908933
transform 1 0 26256 0 1 12913
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_5
timestamp 1626908933
transform 1 0 25920 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_45
timestamp 1626908933
transform 1 0 25920 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_3
timestamp 1626908933
transform 1 0 24192 0 1 13320
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_1
timestamp 1626908933
transform 1 0 24192 0 1 13320
box -38 -49 2726 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_31
timestamp 1626908933
transform 1 0 24192 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_15
timestamp 1626908933
transform 1 0 24192 0 -1 13320
box -38 -49 1670 715
use L1M1_PR  L1M1_PR_1329
timestamp 1626908933
transform 1 0 26832 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1303
timestamp 1626908933
transform 1 0 26640 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_541
timestamp 1626908933
transform 1 0 26832 0 1 12543
box -29 -23 29 23
use L1M1_PR  L1M1_PR_515
timestamp 1626908933
transform 1 0 26640 0 1 12839
box -29 -23 29 23
use L1M1_PR  L1M1_PR_537
timestamp 1626908933
transform 1 0 26736 0 1 13061
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1325
timestamp 1626908933
transform 1 0 26736 0 1 13061
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_170
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_440
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_170
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_440
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_170
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_440
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_181
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_469
timestamp 1626908933
transform 1 0 26600 0 1 13320
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_453
timestamp 1626908933
transform 1 0 26880 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_85
timestamp 1626908933
transform 1 0 26880 0 1 13320
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1242
timestamp 1626908933
transform 1 0 27024 0 1 12543
box -32 -32 32 32
use M1M2_PR  M1M2_PR_474
timestamp 1626908933
transform 1 0 27024 0 1 12543
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1319
timestamp 1626908933
transform 1 0 27408 0 1 12765
box -29 -23 29 23
use L1M1_PR  L1M1_PR_531
timestamp 1626908933
transform 1 0 27408 0 1 12765
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1233
timestamp 1626908933
transform 1 0 27408 0 1 12765
box -32 -32 32 32
use M1M2_PR  M1M2_PR_465
timestamp 1626908933
transform 1 0 27408 0 1 12765
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_355
timestamp 1626908933
transform 1 0 27456 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_96
timestamp 1626908933
transform 1 0 27456 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_457
timestamp 1626908933
transform 1 0 27552 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_89
timestamp 1626908933
transform 1 0 27552 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_738
timestamp 1626908933
transform 1 0 27072 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_169
timestamp 1626908933
transform 1 0 27072 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_14
timestamp 1626908933
transform 1 0 26688 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_54
timestamp 1626908933
transform 1 0 26688 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_133
timestamp 1626908933
transform 1 0 27744 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_763
timestamp 1626908933
transform 1 0 27744 0 -1 13320
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_22
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_310
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_290
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_20
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_290
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_20
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_290
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_20
timestamp 1626908933
transform 1 0 28600 0 1 12654
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_762
timestamp 1626908933
transform 1 0 28800 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_132
timestamp 1626908933
transform 1 0 28800 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_456
timestamp 1626908933
transform 1 0 28608 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_88
timestamp 1626908933
transform 1 0 28608 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_136
timestamp 1626908933
transform 1 0 28896 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_160
timestamp 1626908933
transform 1 0 27840 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_706
timestamp 1626908933
transform 1 0 28896 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_730
timestamp 1626908933
transform 1 0 27840 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_25
timestamp 1626908933
transform 1 0 27456 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_9
timestamp 1626908933
transform 1 0 27456 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_130
timestamp 1626908933
transform 1 0 29184 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_699
timestamp 1626908933
transform 1 0 29184 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_124
timestamp 1626908933
transform 1 0 29088 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_754
timestamp 1626908933
transform 1 0 29088 0 1 13320
box -38 -49 134 715
use M1M2_PR  M1M2_PR_382
timestamp 1626908933
transform 1 0 29616 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_413
timestamp 1626908933
transform 1 0 29712 0 1 12987
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1150
timestamp 1626908933
transform 1 0 29616 0 1 12913
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1181
timestamp 1626908933
transform 1 0 29712 0 1 12987
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_88
timestamp 1626908933
transform 1 0 29568 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_347
timestamp 1626908933
transform 1 0 29568 0 1 13320
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_453
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_165
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_155
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_425
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_155
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_425
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_155
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_425
timestamp 1626908933
transform 1 0 30600 0 1 13320
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_662
timestamp 1626908933
transform 1 0 31296 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_93
timestamp 1626908933
transform 1 0 31296 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_654
timestamp 1626908933
transform 1 0 31680 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_84
timestamp 1626908933
transform 1 0 31680 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_663
timestamp 1626908933
transform 1 0 31296 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_94
timestamp 1626908933
transform 1 0 31296 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_655
timestamp 1626908933
transform 1 0 31680 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_85
timestamp 1626908933
transform 1 0 31680 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_16
timestamp 1626908933
transform 1 0 29664 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_0
timestamp 1626908933
transform 1 0 29664 0 1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_17
timestamp 1626908933
transform 1 0 29664 0 -1 13320
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_1
timestamp 1626908933
transform 1 0 29664 0 -1 13320
box -38 -49 1670 715
use osc_core_VIA4  osc_core_VIA4_294
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_6
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_275
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_5
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_275
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_5
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_275
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_5
timestamp 1626908933
transform 1 0 32600 0 1 12654
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_753
timestamp 1626908933
transform 1 0 32448 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_123
timestamp 1626908933
transform 1 0 32448 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_354
timestamp 1626908933
transform 1 0 32448 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_95
timestamp 1626908933
transform 1 0 32448 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_61
timestamp 1626908933
transform 1 0 32544 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_630
timestamp 1626908933
transform 1 0 32544 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_60
timestamp 1626908933
transform 1 0 32544 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_629
timestamp 1626908933
transform 1 0 32544 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_624
timestamp 1626908933
transform 1 0 32928 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_54
timestamp 1626908933
transform 1 0 32928 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_625
timestamp 1626908933
transform 1 0 32928 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_55
timestamp 1626908933
transform 1 0 32928 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_131
timestamp 1626908933
transform 1 0 33696 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_761
timestamp 1626908933
transform 1 0 33696 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_122
timestamp 1626908933
transform 1 0 33696 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_752
timestamp 1626908933
transform 1 0 33696 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_25
timestamp 1626908933
transform 1 0 34176 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_595
timestamp 1626908933
transform 1 0 34176 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_28
timestamp 1626908933
transform 1 0 33792 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_597
timestamp 1626908933
transform 1 0 33792 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_24
timestamp 1626908933
transform 1 0 34176 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_594
timestamp 1626908933
transform 1 0 34176 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_27
timestamp 1626908933
transform 1 0 33792 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_596
timestamp 1626908933
transform 1 0 33792 0 1 13320
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_410
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_140
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_410
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_140
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_410
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_140
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_149
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_437
timestamp 1626908933
transform 1 0 34600 0 1 13320
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_690
timestamp 1626908933
transform 1 0 35424 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_322
timestamp 1626908933
transform 1 0 35424 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_574
timestamp 1626908933
transform 1 0 35040 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_5
timestamp 1626908933
transform 1 0 35040 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_346
timestamp 1626908933
transform 1 0 34944 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_87
timestamp 1626908933
transform 1 0 34944 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_575
timestamp 1626908933
transform 1 0 34944 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_5
timestamp 1626908933
transform 1 0 34944 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1182
timestamp 1626908933
transform 1 0 35616 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_552
timestamp 1626908933
transform 1 0 35616 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_30
timestamp 1626908933
transform 1 0 288 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_5
timestamp 1626908933
transform 1 0 288 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1415
timestamp 1626908933
transform 1 0 144 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_647
timestamp 1626908933
transform 1 0 144 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1139
timestamp 1626908933
transform 1 0 624 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_351
timestamp 1626908933
transform 1 0 624 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1465
timestamp 1626908933
transform 1 0 432 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_677
timestamp 1626908933
transform 1 0 432 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1198
timestamp 1626908933
transform 1 0 720 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_410
timestamp 1626908933
transform 1 0 720 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1259
timestamp 1626908933
transform 1 0 528 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_471
timestamp 1626908933
transform 1 0 528 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1164
timestamp 1626908933
transform 1 0 528 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_396
timestamp 1626908933
transform 1 0 528 0 1 13653
box -32 -32 32 32
use M2M3_PR  M2M3_PR_85
timestamp 1626908933
transform 1 0 528 0 1 13701
box -33 -37 33 37
use M2M3_PR  M2M3_PR_26
timestamp 1626908933
transform 1 0 528 0 1 13701
box -33 -37 33 37
use osc_core_VIA7  osc_core_VIA7_394
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_124
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_394
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_124
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_394
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_124
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_133
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_421
timestamp 1626908933
transform 1 0 600 0 1 13986
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_323
timestamp 1626908933
transform 1 0 672 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_691
timestamp 1626908933
transform 1 0 672 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_97
timestamp 1626908933
transform -1 0 1344 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_42
timestamp 1626908933
transform -1 0 1344 0 -1 14652
box -38 -49 518 715
use M1M2_PR  M1M2_PR_290
timestamp 1626908933
transform 1 0 1008 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1058
timestamp 1626908933
transform 1 0 1008 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_354
timestamp 1626908933
transform 1 0 1008 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1142
timestamp 1626908933
transform 1 0 1008 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_332
timestamp 1626908933
transform 1 0 1104 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1100
timestamp 1626908933
transform 1 0 1104 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_285
timestamp 1626908933
transform 1 0 1296 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1053
timestamp 1626908933
transform 1 0 1296 0 1 13431
box -32 -32 32 32
use L1M1_PR  L1M1_PR_193
timestamp 1626908933
transform 1 0 1200 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_981
timestamp 1626908933
transform 1 0 1200 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_324
timestamp 1626908933
transform 1 0 1344 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_692
timestamp 1626908933
transform 1 0 1344 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_283
timestamp 1626908933
transform 1 0 1776 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1051
timestamp 1626908933
transform 1 0 1776 0 1 13431
box -32 -32 32 32
use L1M1_PR  L1M1_PR_345
timestamp 1626908933
transform 1 0 1776 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1133
timestamp 1626908933
transform 1 0 1776 0 1 13431
box -29 -23 29 23
use M1M2_PR  M1M2_PR_149
timestamp 1626908933
transform 1 0 1488 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_917
timestamp 1626908933
transform 1 0 1488 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_386
timestamp 1626908933
transform 1 0 1680 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1154
timestamp 1626908933
transform 1 0 1680 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_459
timestamp 1626908933
transform 1 0 1680 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1247
timestamp 1626908933
transform 1 0 1680 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1412
timestamp 1626908933
transform 1 0 1488 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_644
timestamp 1626908933
transform 1 0 1488 0 1 13875
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1463
timestamp 1626908933
transform 1 0 1488 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_675
timestamp 1626908933
transform 1 0 1488 0 1 13875
box -29 -23 29 23
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_47
timestamp 1626908933
transform 1 0 1536 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_22
timestamp 1626908933
transform 1 0 1536 0 -1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1210
timestamp 1626908933
transform 1 0 1968 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_422
timestamp 1626908933
transform 1 0 1968 0 1 13875
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1183
timestamp 1626908933
transform 1 0 1920 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_553
timestamp 1626908933
transform 1 0 1920 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1039
timestamp 1626908933
transform 1 0 2064 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_271
timestamp 1626908933
transform 1 0 2064 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1114
timestamp 1626908933
transform 1 0 2256 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_346
timestamp 1626908933
transform 1 0 2256 0 1 13875
box -32 -32 32 32
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_44
timestamp 1626908933
transform 1 0 2016 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_19
timestamp 1626908933
transform 1 0 2016 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_268
timestamp 1626908933
transform 1 0 2448 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1036
timestamp 1626908933
transform 1 0 2448 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_114
timestamp 1626908933
transform 1 0 2544 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_329
timestamp 1626908933
transform 1 0 2352 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_902
timestamp 1626908933
transform 1 0 2544 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1117
timestamp 1626908933
transform 1 0 2352 0 1 13579
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_86
timestamp 1626908933
transform 1 0 2496 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_345
timestamp 1626908933
transform 1 0 2496 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_554
timestamp 1626908933
transform 1 0 2400 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1184
timestamp 1626908933
transform 1 0 2400 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_751
timestamp 1626908933
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_121
timestamp 1626908933
transform 1 0 2592 0 -1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1120
timestamp 1626908933
transform 1 0 2736 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_332
timestamp 1626908933
transform 1 0 2736 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1108
timestamp 1626908933
transform 1 0 2688 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_539
timestamp 1626908933
transform 1 0 2688 0 -1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_111
timestamp 1626908933
transform 1 0 2928 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_899
timestamp 1626908933
transform 1 0 2928 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1089
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_321
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -32 -32 32 32
use M3M4_PR  M3M4_PR_38
timestamp 1626908933
transform 1 0 3552 0 1 13701
box -38 -33 38 33
use M3M4_PR  M3M4_PR_17
timestamp 1626908933
transform 1 0 3552 0 1 13701
box -38 -33 38 33
use L1M1_PR  L1M1_PR_1182
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_394
timestamp 1626908933
transform 1 0 3504 0 1 13653
box -29 -23 29 23
use M2M3_PR  M2M3_PR_77
timestamp 1626908933
transform 1 0 3600 0 1 13701
box -33 -37 33 37
use M2M3_PR  M2M3_PR_18
timestamp 1626908933
transform 1 0 3600 0 1 13701
box -33 -37 33 37
use L1M1_PR  L1M1_PR_972
timestamp 1626908933
transform 1 0 3600 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_184
timestamp 1626908933
transform 1 0 3600 0 1 13727
box -29 -23 29 23
use M1M2_PR  M1M2_PR_915
timestamp 1626908933
transform 1 0 3600 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_147
timestamp 1626908933
transform 1 0 3600 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_27
timestamp 1626908933
transform 1 0 3072 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_2
timestamp 1626908933
transform 1 0 3072 0 -1 14652
box -38 -49 1670 715
use osc_core_VIA4  osc_core_VIA4_405
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_117
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -142 200 178
use L1M1_PR  L1M1_PR_896
timestamp 1626908933
transform 1 0 4368 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_108
timestamp 1626908933
transform 1 0 4368 0 1 13653
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_379
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_109
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_379
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_109
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_379
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_109
timestamp 1626908933
transform 1 0 4600 0 1 13986
box -200 -49 200 49
use M1M2_PR  M1M2_PR_86
timestamp 1626908933
transform 1 0 4944 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_854
timestamp 1626908933
transform 1 0 4944 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_555
timestamp 1626908933
transform 1 0 4704 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1185
timestamp 1626908933
transform 1 0 4704 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_84
timestamp 1626908933
transform -1 0 5280 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_29
timestamp 1626908933
transform -1 0 5280 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_750
timestamp 1626908933
transform 1 0 5280 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_120
timestamp 1626908933
transform 1 0 5280 0 -1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1129
timestamp 1626908933
transform 1 0 5232 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_341
timestamp 1626908933
transform 1 0 5232 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1047
timestamp 1626908933
transform 1 0 5232 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_279
timestamp 1626908933
transform 1 0 5232 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_884
timestamp 1626908933
transform 1 0 5424 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_96
timestamp 1626908933
transform 1 0 5424 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1082
timestamp 1626908933
transform 1 0 5376 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_513
timestamp 1626908933
transform 1 0 5376 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_264
timestamp 1626908933
transform 1 0 6000 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1032
timestamp 1626908933
transform 1 0 6000 0 1 13431
box -32 -32 32 32
use L1M1_PR  L1M1_PR_325
timestamp 1626908933
transform 1 0 6000 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1113
timestamp 1626908933
transform 1 0 6000 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_28
timestamp 1626908933
transform 1 0 5760 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_108
timestamp 1626908933
transform 1 0 5760 0 -1 14652
box -38 -49 902 715
use M1M2_PR  M1M2_PR_32
timestamp 1626908933
transform 1 0 6192 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_800
timestamp 1626908933
transform 1 0 6192 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_37
timestamp 1626908933
transform 1 0 6192 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_825
timestamp 1626908933
transform 1 0 6192 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_737
timestamp 1626908933
transform 1 0 6864 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1505
timestamp 1626908933
transform 1 0 6864 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_762
timestamp 1626908933
transform 1 0 6864 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1550
timestamp 1626908933
transform 1 0 6864 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_31
timestamp 1626908933
transform 1 0 6624 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_111
timestamp 1626908933
transform 1 0 6624 0 -1 14652
box -38 -49 902 715
use M1M2_PR  M1M2_PR_27
timestamp 1626908933
transform 1 0 7152 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_795
timestamp 1626908933
transform 1 0 7152 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_29
timestamp 1626908933
transform 1 0 7152 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_817
timestamp 1626908933
transform 1 0 7152 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_85
timestamp 1626908933
transform 1 0 7488 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_344
timestamp 1626908933
transform 1 0 7488 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_112
timestamp 1626908933
transform 1 0 8112 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_880
timestamp 1626908933
transform 1 0 8112 0 1 13727
box -32 -32 32 32
use L1M1_PR  L1M1_PR_131
timestamp 1626908933
transform 1 0 8112 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_919
timestamp 1626908933
transform 1 0 8112 0 1 13727
box -29 -23 29 23
use M2M3_PR  M2M3_PR_10
timestamp 1626908933
transform 1 0 8112 0 1 13701
box -33 -37 33 37
use M2M3_PR  M2M3_PR_69
timestamp 1626908933
transform 1 0 8112 0 1 13701
box -33 -37 33 37
use M3M4_PR  M3M4_PR_9
timestamp 1626908933
transform 1 0 8112 0 1 13701
box -38 -33 38 33
use M3M4_PR  M3M4_PR_30
timestamp 1626908933
transform 1 0 8112 0 1 13701
box -38 -33 38 33
use M1M2_PR  M1M2_PR_316
timestamp 1626908933
transform 1 0 8304 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1084
timestamp 1626908933
transform 1 0 8304 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_387
timestamp 1626908933
transform 1 0 8304 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1175
timestamp 1626908933
transform 1 0 8304 0 1 13653
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_101
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_389
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -142 200 178
use L1M1_PR  L1M1_PR_954
timestamp 1626908933
transform 1 0 8976 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_166
timestamp 1626908933
transform 1 0 8976 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_900
timestamp 1626908933
transform 1 0 8976 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_132
timestamp 1626908933
transform 1 0 8976 0 1 13653
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_364
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_94
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_364
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_94
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_364
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_94
timestamp 1626908933
transform 1 0 8600 0 1 13986
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_556
timestamp 1626908933
transform 1 0 9216 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1186
timestamp 1626908933
transform 1 0 9216 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_49
timestamp 1626908933
transform -1 0 10176 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_129
timestamp 1626908933
transform -1 0 10176 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_47
timestamp 1626908933
transform 1 0 7584 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_22
timestamp 1626908933
transform 1 0 7584 0 -1 14652
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_22
timestamp 1626908933
transform 1 0 9840 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_790
timestamp 1626908933
transform 1 0 9840 0 1 13431
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_325
timestamp 1626908933
transform 1 0 10176 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_693
timestamp 1626908933
transform 1 0 10176 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_682
timestamp 1626908933
transform 1 0 10512 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1450
timestamp 1626908933
transform 1 0 10512 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_716
timestamp 1626908933
transform 1 0 10512 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1504
timestamp 1626908933
transform 1 0 10512 0 1 13653
box -29 -23 29 23
use M2M3_PR  M2M3_PR_52
timestamp 1626908933
transform 1 0 10512 0 1 13701
box -33 -37 33 37
use M2M3_PR  M2M3_PR_111
timestamp 1626908933
transform 1 0 10512 0 1 13701
box -33 -37 33 37
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_50
timestamp 1626908933
transform 1 0 10368 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_130
timestamp 1626908933
transform 1 0 10368 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_133
timestamp 1626908933
transform 1 0 11424 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_53
timestamp 1626908933
transform 1 0 11424 0 -1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_694
timestamp 1626908933
transform 1 0 11232 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_326
timestamp 1626908933
transform 1 0 11232 0 -1 14652
box -38 -49 230 715
use L1M1_PR  L1M1_PR_949
timestamp 1626908933
transform 1 0 10800 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_161
timestamp 1626908933
transform 1 0 10800 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_677
timestamp 1626908933
transform 1 0 11760 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1445
timestamp 1626908933
transform 1 0 11760 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_710
timestamp 1626908933
transform 1 0 11760 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1498
timestamp 1626908933
transform 1 0 11760 0 1 13653
box -29 -23 29 23
use M2M3_PR  M2M3_PR_51
timestamp 1626908933
transform 1 0 11760 0 1 13701
box -33 -37 33 37
use M2M3_PR  M2M3_PR_110
timestamp 1626908933
transform 1 0 11760 0 1 13701
box -33 -37 33 37
use M1M2_PR  M1M2_PR_72
timestamp 1626908933
transform 1 0 12144 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_840
timestamp 1626908933
transform 1 0 12144 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_82
timestamp 1626908933
transform 1 0 12144 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_870
timestamp 1626908933
transform 1 0 12144 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_327
timestamp 1626908933
transform 1 0 12288 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_695
timestamp 1626908933
transform 1 0 12288 0 -1 14652
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_79
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_349
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_79
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_349
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_79
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_349
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_85
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_373
timestamp 1626908933
transform 1 0 12600 0 1 13986
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_394
timestamp 1626908933
transform 1 0 12768 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_963
timestamp 1626908933
transform 1 0 12768 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_84
timestamp 1626908933
transform 1 0 12576 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_452
timestamp 1626908933
transform 1 0 12576 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_84
timestamp 1626908933
transform 1 0 12480 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_343
timestamp 1626908933
transform 1 0 12480 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_310
timestamp 1626908933
transform 1 0 13680 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1078
timestamp 1626908933
transform 1 0 13680 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_382
timestamp 1626908933
transform 1 0 13680 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1170
timestamp 1626908933
transform 1 0 13680 0 1 13653
box -29 -23 29 23
use osc_core_VIA0  osc_core_VIA0_3
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_8
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_3
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_8
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -33 96 33
use osc_core_VIA2  osc_core_VIA2_3
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_8
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_3
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_8
timestamp 1626908933
transform 1 0 14116 0 1 13502
box -97 -28 96 28
use M1M2_PR  M1M2_PR_13
timestamp 1626908933
transform 1 0 14640 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_781
timestamp 1626908933
transform 1 0 14640 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_8
timestamp 1626908933
transform 1 0 14640 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_796
timestamp 1626908933
transform 1 0 14640 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_83
timestamp 1626908933
transform 1 0 14784 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_451
timestamp 1626908933
transform 1 0 14784 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_407
timestamp 1626908933
transform 1 0 14976 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_977
timestamp 1626908933
transform 1 0 14976 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_32
timestamp 1626908933
transform 1 0 13152 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_7
timestamp 1626908933
transform 1 0 13152 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_343
timestamp 1626908933
transform 1 0 15840 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_912
timestamp 1626908933
transform 1 0 15840 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_119
timestamp 1626908933
transform 1 0 15744 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_749
timestamp 1626908933
transform 1 0 15744 0 -1 14652
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_64
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_334
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_64
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_334
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_64
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_334
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_69
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_357
timestamp 1626908933
transform 1 0 16600 0 1 13986
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_378
timestamp 1626908933
transform 1 0 16224 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_948
timestamp 1626908933
transform 1 0 16224 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_342
timestamp 1626908933
transform 1 0 17376 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_83
timestamp 1626908933
transform 1 0 17376 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_888
timestamp 1626908933
transform 1 0 16992 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_319
timestamp 1626908933
transform 1 0 16992 0 -1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_814
timestamp 1626908933
transform 1 0 18000 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_46
timestamp 1626908933
transform 1 0 18000 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_42
timestamp 1626908933
transform 1 0 17472 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_17
timestamp 1626908933
transform 1 0 17472 0 -1 14652
box -38 -49 1670 715
use L1M1_PR  L1M1_PR_839
timestamp 1626908933
transform 1 0 18000 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_51
timestamp 1626908933
transform 1 0 18000 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1410
timestamp 1626908933
transform 1 0 18288 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_622
timestamp 1626908933
transform 1 0 18288 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1315
timestamp 1626908933
transform 1 0 18288 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_547
timestamp 1626908933
transform 1 0 18288 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_101
timestamp 1626908933
transform 1 0 19056 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_869
timestamp 1626908933
transform 1 0 19056 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_117
timestamp 1626908933
transform 1 0 18960 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_905
timestamp 1626908933
transform 1 0 18960 0 1 13653
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_82
timestamp 1626908933
transform 1 0 19104 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_450
timestamp 1626908933
transform 1 0 19104 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_118
timestamp 1626908933
transform 1 0 19296 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_748
timestamp 1626908933
transform 1 0 19296 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_313
timestamp 1626908933
transform 1 0 19392 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_883
timestamp 1626908933
transform 1 0 19392 0 -1 14652
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_341
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_53
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_319
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_49
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_319
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_49
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_319
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_49
timestamp 1626908933
transform 1 0 20600 0 1 13986
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_747
timestamp 1626908933
transform 1 0 20160 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_117
timestamp 1626908933
transform 1 0 20160 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_266
timestamp 1626908933
transform 1 0 20256 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_835
timestamp 1626908933
transform 1 0 20256 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_857
timestamp 1626908933
transform 1 0 20640 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_287
timestamp 1626908933
transform 1 0 20640 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_341
timestamp 1626908933
transform 1 0 21408 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_82
timestamp 1626908933
transform 1 0 21408 0 -1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1417
timestamp 1626908933
transform 1 0 21936 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_629
timestamp 1626908933
transform 1 0 21936 0 1 13653
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1321
timestamp 1626908933
transform 1 0 21936 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_553
timestamp 1626908933
transform 1 0 21936 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2
timestamp 1626908933
transform 1 0 22320 0 1 13505
box -32 -32 32 32
use M1M2_PR  M1M2_PR_770
timestamp 1626908933
transform 1 0 22320 0 1 13505
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1
timestamp 1626908933
transform 1 0 22416 0 1 13505
box -29 -23 29 23
use L1M1_PR  L1M1_PR_789
timestamp 1626908933
transform 1 0 22416 0 1 13505
box -29 -23 29 23
use M1M2_PR  M1M2_PR_39
timestamp 1626908933
transform 1 0 22992 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_807
timestamp 1626908933
transform 1 0 22992 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_42
timestamp 1626908933
transform 1 0 22992 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_830
timestamp 1626908933
transform 1 0 22992 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_500
timestamp 1626908933
transform 1 0 23472 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1288
timestamp 1626908933
transform 1 0 23472 0 1 13727
box -29 -23 29 23
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_17
timestamp 1626908933
transform 1 0 23136 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_57
timestamp 1626908933
transform 1 0 23136 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_37
timestamp 1626908933
transform 1 0 21504 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_12
timestamp 1626908933
transform 1 0 21504 0 -1 14652
box -38 -49 1670 715
use L1M1_PR  L1M1_PR_441
timestamp 1626908933
transform 1 0 23856 0 1 13431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1229
timestamp 1626908933
transform 1 0 23856 0 1 13431
box -29 -23 29 23
use M1M2_PR  M1M2_PR_366
timestamp 1626908933
transform 1 0 23664 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1134
timestamp 1626908933
transform 1 0 23664 0 1 13579
box -32 -32 32 32
use L1M1_PR  L1M1_PR_439
timestamp 1626908933
transform 1 0 23664 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1227
timestamp 1626908933
transform 1 0 23664 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_438
timestamp 1626908933
transform 1 0 23760 0 1 13579
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1226
timestamp 1626908933
transform 1 0 23760 0 1 13579
box -29 -23 29 23
use M1M2_PR  M1M2_PR_364
timestamp 1626908933
transform 1 0 23856 0 1 13579
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1132
timestamp 1626908933
transform 1 0 23856 0 1 13579
box -32 -32 32 32
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_0
timestamp 1626908933
transform 1 0 23904 0 -1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__conb_1  sky130_fd_sc_hs__conb_1_1
timestamp 1626908933
transform 1 0 23904 0 -1 14652
box -38 -49 326 715
use M1M2_PR  M1M2_PR_1138
timestamp 1626908933
transform 1 0 24144 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_370
timestamp 1626908933
transform 1 0 24144 0 1 13431
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1136
timestamp 1626908933
transform 1 0 24048 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_368
timestamp 1626908933
transform 1 0 24048 0 1 13653
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1228
timestamp 1626908933
transform 1 0 24048 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_440
timestamp 1626908933
transform 1 0 24048 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1293
timestamp 1626908933
transform 1 0 24240 0 1 13727
box -29 -23 29 23
use L1M1_PR  L1M1_PR_505
timestamp 1626908933
transform 1 0 24240 0 1 13727
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1216
timestamp 1626908933
transform 1 0 24144 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_448
timestamp 1626908933
transform 1 0 24144 0 1 13727
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_325
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_37
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1268
timestamp 1626908933
transform 1 0 24624 0 1 13653
box -29 -23 29 23
use L1M1_PR  L1M1_PR_480
timestamp 1626908933
transform 1 0 24624 0 1 13653
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_304
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_34
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_304
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_34
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_304
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_34
timestamp 1626908933
transform 1 0 24600 0 1 13986
box -200 -49 200 49
use M1M2_PR  M1M2_PR_406
timestamp 1626908933
transform 1 0 24912 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1174
timestamp 1626908933
transform 1 0 24912 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1209
timestamp 1626908933
transform 1 0 25488 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_441
timestamp 1626908933
transform 1 0 25488 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_2
timestamp 1626908933
transform 1 0 24192 0 -1 14652
box -38 -49 2726 715
use sky130_fd_sc_hs__dfrtp_4  sky130_fd_sc_hs__dfrtp_4_0
timestamp 1626908933
transform 1 0 24192 0 -1 14652
box -38 -49 2726 715
use M1M2_PR  M1M2_PR_363
timestamp 1626908933
transform 1 0 26640 0 1 13875
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1131
timestamp 1626908933
transform 1 0 26640 0 1 13875
box -32 -32 32 32
use L1M1_PR  L1M1_PR_435
timestamp 1626908933
transform 1 0 26448 0 1 13875
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1223
timestamp 1626908933
transform 1 0 26448 0 1 13875
box -29 -23 29 23
use M1M2_PR  M1M2_PR_373
timestamp 1626908933
transform 1 0 27216 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1141
timestamp 1626908933
transform 1 0 27216 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_0
timestamp 1626908933
transform 1 0 26880 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_2
timestamp 1626908933
transform 1 0 26880 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_81
timestamp 1626908933
transform 1 0 27360 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_340
timestamp 1626908933
transform 1 0 27360 0 -1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_426
timestamp 1626908933
transform 1 0 29040 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1194
timestamp 1626908933
transform 1 0 29040 0 1 13653
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_19
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_289
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_19
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_289
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_19
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_289
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_21
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_309
timestamp 1626908933
transform 1 0 28600 0 1 13986
box -200 -142 200 178
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_24
timestamp 1626908933
transform 1 0 27456 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_8
timestamp 1626908933
transform 1 0 27456 0 -1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_81
timestamp 1626908933
transform 1 0 29088 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_449
timestamp 1626908933
transform 1 0 29088 0 -1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_411
timestamp 1626908933
transform 1 0 29712 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_412
timestamp 1626908933
transform 1 0 29808 0 1 13727
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1179
timestamp 1626908933
transform 1 0 29712 0 1 13653
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1180
timestamp 1626908933
transform 1 0 29808 0 1 13727
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_27
timestamp 1626908933
transform 1 0 29664 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_7
timestamp 1626908933
transform 1 0 29664 0 -1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_129
timestamp 1626908933
transform 1 0 29280 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_698
timestamp 1626908933
transform 1 0 29280 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_339
timestamp 1626908933
transform 1 0 30144 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_80
timestamp 1626908933
transform 1 0 30144 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_746
timestamp 1626908933
transform 1 0 30240 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_116
timestamp 1626908933
transform 1 0 30240 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_683
timestamp 1626908933
transform 1 0 30336 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_113
timestamp 1626908933
transform 1 0 30336 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_448
timestamp 1626908933
transform 1 0 31104 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_80
timestamp 1626908933
transform 1 0 31104 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_661
timestamp 1626908933
transform 1 0 31296 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_92
timestamp 1626908933
transform 1 0 31296 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_653
timestamp 1626908933
transform 1 0 31680 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_83
timestamp 1626908933
transform 1 0 31680 0 -1 14652
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_293
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_5
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_274
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_4
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_274
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_4
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_274
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_4
timestamp 1626908933
transform 1 0 32600 0 1 13986
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_338
timestamp 1626908933
transform 1 0 32448 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_79
timestamp 1626908933
transform 1 0 32448 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_59
timestamp 1626908933
transform 1 0 32544 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_628
timestamp 1626908933
transform 1 0 32544 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_623
timestamp 1626908933
transform 1 0 32928 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_53
timestamp 1626908933
transform 1 0 32928 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_745
timestamp 1626908933
transform 1 0 33696 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_115
timestamp 1626908933
transform 1 0 33696 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_595
timestamp 1626908933
transform 1 0 33792 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_26
timestamp 1626908933
transform 1 0 33792 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_593
timestamp 1626908933
transform 1 0 34176 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_23
timestamp 1626908933
transform 1 0 34176 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_4
timestamp 1626908933
transform 1 0 34944 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_574
timestamp 1626908933
transform 1 0 34944 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_337
timestamp 1626908933
transform 1 0 288 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_78
timestamp 1626908933
transform 1 0 288 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1419
timestamp 1626908933
transform 1 0 48 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_651
timestamp 1626908933
transform 1 0 48 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1416
timestamp 1626908933
transform 1 0 48 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_648
timestamp 1626908933
transform 1 0 48 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1264
timestamp 1626908933
transform 1 0 432 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_476
timestamp 1626908933
transform 1 0 432 0 1 14319
box -29 -23 29 23
use M2M3_PR  M2M3_PR_84
timestamp 1626908933
transform 1 0 528 0 1 14311
box -33 -37 33 37
use M2M3_PR  M2M3_PR_25
timestamp 1626908933
transform 1 0 528 0 1 14311
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1163
timestamp 1626908933
transform 1 0 528 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_395
timestamp 1626908933
transform 1 0 528 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1466
timestamp 1626908933
transform 1 0 336 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_678
timestamp 1626908933
transform 1 0 336 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1145
timestamp 1626908933
transform 1 0 528 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_357
timestamp 1626908933
transform 1 0 528 0 1 14541
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1187
timestamp 1626908933
transform 1 0 576 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_557
timestamp 1626908933
transform 1 0 576 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_696
timestamp 1626908933
transform 1 0 384 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_328
timestamp 1626908933
transform 1 0 384 0 1 14652
box -38 -49 230 715
use L1M1_PR  L1M1_PR_356
timestamp 1626908933
transform 1 0 624 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_417
timestamp 1626908933
transform 1 0 624 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1144
timestamp 1626908933
transform 1 0 624 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1205
timestamp 1626908933
transform 1 0 624 0 1 14393
box -29 -23 29 23
use M1M2_PR  M1M2_PR_292
timestamp 1626908933
transform 1 0 624 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1060
timestamp 1626908933
transform 1 0 624 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_92
timestamp 1626908933
transform 1 0 672 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_37
timestamp 1626908933
transform 1 0 672 0 1 14652
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1057
timestamp 1626908933
transform 1 0 1008 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_289
timestamp 1626908933
transform 1 0 1008 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_986
timestamp 1626908933
transform 1 0 1008 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_198
timestamp 1626908933
transform 1 0 1008 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_923
timestamp 1626908933
transform 1 0 1008 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_155
timestamp 1626908933
transform 1 0 1008 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1150
timestamp 1626908933
transform 1 0 1200 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_362
timestamp 1626908933
transform 1 0 1200 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1107
timestamp 1626908933
transform 1 0 1104 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_339
timestamp 1626908933
transform 1 0 1104 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_294
timestamp 1626908933
transform 1 0 1296 0 1 14467
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1062
timestamp 1626908933
transform 1 0 1296 0 1 14467
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_96
timestamp 1626908933
transform 1 0 1152 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_41
timestamp 1626908933
transform 1 0 1152 0 1 14652
box -38 -49 518 715
use M2M3_PR  M2M3_PR_83
timestamp 1626908933
transform 1 0 1680 0 1 14311
box -33 -37 33 37
use M2M3_PR  M2M3_PR_24
timestamp 1626908933
transform 1 0 1680 0 1 14311
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1153
timestamp 1626908933
transform 1 0 1680 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_385
timestamp 1626908933
transform 1 0 1680 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1246
timestamp 1626908933
transform 1 0 1680 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_458
timestamp 1626908933
transform 1 0 1680 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1411
timestamp 1626908933
transform 1 0 1488 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_643
timestamp 1626908933
transform 1 0 1488 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1462
timestamp 1626908933
transform 1 0 1584 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_674
timestamp 1626908933
transform 1 0 1584 0 1 14393
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_329
timestamp 1626908933
transform 1 0 1632 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_697
timestamp 1626908933
transform 1 0 1632 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1122
timestamp 1626908933
transform 1 0 1872 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_354
timestamp 1626908933
transform 1 0 1872 0 1 14763
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1216
timestamp 1626908933
transform 1 0 1872 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1146
timestamp 1626908933
transform 1 0 1776 0 1 14467
box -29 -23 29 23
use L1M1_PR  L1M1_PR_428
timestamp 1626908933
transform 1 0 1872 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_358
timestamp 1626908933
transform 1 0 1776 0 1 14467
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1123
timestamp 1626908933
transform 1 0 1872 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_355
timestamp 1626908933
transform 1 0 1872 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_39
timestamp 1626908933
transform -1 0 2304 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_94
timestamp 1626908933
transform -1 0 2304 0 1 14652
box -38 -49 518 715
use L1M1_PR  L1M1_PR_328
timestamp 1626908933
transform 1 0 2352 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1116
timestamp 1626908933
transform 1 0 2352 0 1 14097
box -29 -23 29 23
use M1M2_PR  M1M2_PR_267
timestamp 1626908933
transform 1 0 2448 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1035
timestamp 1626908933
transform 1 0 2448 0 1 14097
box -32 -32 32 32
use L1M1_PR  L1M1_PR_681
timestamp 1626908933
transform 1 0 1968 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1469
timestamp 1626908933
transform 1 0 1968 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_454
timestamp 1626908933
transform 1 0 2160 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1242
timestamp 1626908933
transform 1 0 2160 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_420
timestamp 1626908933
transform 1 0 2352 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1208
timestamp 1626908933
transform 1 0 2352 0 1 14393
box -29 -23 29 23
use M1M2_PR  M1M2_PR_345
timestamp 1626908933
transform 1 0 2256 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1113
timestamp 1626908933
transform 1 0 2256 0 1 14393
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1468
timestamp 1626908933
transform 1 0 1968 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_680
timestamp 1626908933
transform 1 0 1968 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1418
timestamp 1626908933
transform 1 0 2160 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_650
timestamp 1626908933
transform 1 0 2160 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1331
timestamp 1626908933
transform 1 0 2352 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_563
timestamp 1626908933
transform 1 0 2352 0 1 14541
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_529
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_259
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_529
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_259
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_529
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_259
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_276
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_564
timestamp 1626908933
transform 1 0 2600 0 1 14652
box -200 -142 200 178
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_45
timestamp 1626908933
transform 1 0 2304 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__a21oi_1  sky130_fd_sc_hs__a21oi_1_20
timestamp 1626908933
transform 1 0 2304 0 1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_424
timestamp 1626908933
transform 1 0 2736 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1212
timestamp 1626908933
transform 1 0 2736 0 1 14763
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_5
timestamp 1626908933
transform 1 0 2688 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_14
timestamp 1626908933
transform 1 0 2688 0 1 14652
box -38 -49 422 715
use M3M4_PR  M3M4_PR_16
timestamp 1626908933
transform 1 0 3552 0 1 14189
box -38 -33 38 33
use M3M4_PR  M3M4_PR_37
timestamp 1626908933
transform 1 0 3552 0 1 14189
box -38 -33 38 33
use M1M2_PR  M1M2_PR_320
timestamp 1626908933
transform 1 0 3504 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1088
timestamp 1626908933
transform 1 0 3504 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_393
timestamp 1626908933
transform 1 0 3504 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1181
timestamp 1626908933
transform 1 0 3504 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_145
timestamp 1626908933
transform 1 0 3696 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_913
timestamp 1626908933
transform 1 0 3696 0 1 14245
box -32 -32 32 32
use L1M1_PR  L1M1_PR_182
timestamp 1626908933
transform 1 0 3696 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_970
timestamp 1626908933
transform 1 0 3696 0 1 14245
box -29 -23 29 23
use M2M3_PR  M2M3_PR_16
timestamp 1626908933
transform 1 0 3696 0 1 14189
box -33 -37 33 37
use M2M3_PR  M2M3_PR_75
timestamp 1626908933
transform 1 0 3696 0 1 14189
box -33 -37 33 37
use L1M1_PR  L1M1_PR_390
timestamp 1626908933
transform 1 0 3888 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1178
timestamp 1626908933
transform 1 0 3888 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_560
timestamp 1626908933
transform 1 0 4080 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1328
timestamp 1626908933
transform 1 0 4080 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_26
timestamp 1626908933
transform 1 0 3072 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_1
timestamp 1626908933
transform 1 0 3072 0 1 14652
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_91
timestamp 1626908933
transform 1 0 4560 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_859
timestamp 1626908933
transform 1 0 4560 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_105
timestamp 1626908933
transform 1 0 4560 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_893
timestamp 1626908933
transform 1 0 4560 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_90
timestamp 1626908933
transform 1 0 4560 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_858
timestamp 1626908933
transform 1 0 4560 0 1 14837
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1188
timestamp 1626908933
transform 1 0 4896 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_558
timestamp 1626908933
transform 1 0 4896 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_336
timestamp 1626908933
transform 1 0 4992 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_77
timestamp 1626908933
transform 1 0 4992 0 1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_889
timestamp 1626908933
transform 1 0 4944 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_101
timestamp 1626908933
transform 1 0 4944 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_853
timestamp 1626908933
transform 1 0 4944 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_85
timestamp 1626908933
transform 1 0 4944 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_698
timestamp 1626908933
transform 1 0 4704 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_330
timestamp 1626908933
transform 1 0 4704 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_85
timestamp 1626908933
transform 1 0 5088 0 1 14652
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_30
timestamp 1626908933
transform 1 0 5088 0 1 14652
box -38 -49 518 715
use M1M2_PR  M1M2_PR_281
timestamp 1626908933
transform 1 0 5136 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1049
timestamp 1626908933
transform 1 0 5136 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_342
timestamp 1626908933
transform 1 0 5136 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1130
timestamp 1626908933
transform 1 0 5136 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_331
timestamp 1626908933
transform 1 0 5568 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_699
timestamp 1626908933
transform 1 0 5568 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_742
timestamp 1626908933
transform 1 0 6000 0 1 14393
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1510
timestamp 1626908933
transform 1 0 6000 0 1 14393
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_559
timestamp 1626908933
transform 1 0 5760 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1189
timestamp 1626908933
transform 1 0 5760 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_29
timestamp 1626908933
transform 1 0 5856 0 1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_109
timestamp 1626908933
transform 1 0 5856 0 1 14652
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1555
timestamp 1626908933
transform 1 0 6096 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_767
timestamp 1626908933
transform 1 0 6096 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_822
timestamp 1626908933
transform 1 0 6288 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_34
timestamp 1626908933
transform 1 0 6288 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_799
timestamp 1626908933
transform 1 0 6288 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_31
timestamp 1626908933
transform 1 0 6288 0 1 14319
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_548
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_260
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_514
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_244
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_514
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_244
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_514
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_244
timestamp 1626908933
transform 1 0 6600 0 1 14652
box -200 -49 200 49
use M1M2_PR  M1M2_PR_736
timestamp 1626908933
transform 1 0 6864 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1504
timestamp 1626908933
transform 1 0 6864 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_763
timestamp 1626908933
transform 1 0 6768 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1551
timestamp 1626908933
transform 1 0 6768 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_114
timestamp 1626908933
transform 1 0 6720 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_744
timestamp 1626908933
transform 1 0 6720 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_501
timestamp 1626908933
transform 1 0 6816 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1071
timestamp 1626908933
transform 1 0 6816 0 1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_26
timestamp 1626908933
transform 1 0 7152 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_794
timestamp 1626908933
transform 1 0 7152 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_28
timestamp 1626908933
transform 1 0 7152 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_816
timestamp 1626908933
transform 1 0 7152 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_918
timestamp 1626908933
transform 1 0 8112 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_130
timestamp 1626908933
transform 1 0 8112 0 1 14245
box -29 -23 29 23
use M1M2_PR  M1M2_PR_879
timestamp 1626908933
transform 1 0 8112 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_111
timestamp 1626908933
transform 1 0 8112 0 1 14245
box -32 -32 32 32
use M3M4_PR  M3M4_PR_29
timestamp 1626908933
transform 1 0 8112 0 1 14311
box -38 -33 38 33
use M3M4_PR  M3M4_PR_8
timestamp 1626908933
transform 1 0 8112 0 1 14311
box -38 -33 38 33
use M2M3_PR  M2M3_PR_68
timestamp 1626908933
transform 1 0 8112 0 1 14311
box -33 -37 33 37
use M2M3_PR  M2M3_PR_9
timestamp 1626908933
transform 1 0 8112 0 1 14311
box -33 -37 33 37
use L1M1_PR  L1M1_PR_1177
timestamp 1626908933
transform 1 0 8016 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_389
timestamp 1626908933
transform 1 0 8016 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_315
timestamp 1626908933
transform 1 0 8304 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1083
timestamp 1626908933
transform 1 0 8304 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_131
timestamp 1626908933
transform 1 0 8976 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_899
timestamp 1626908933
transform 1 0 8976 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_165
timestamp 1626908933
transform 1 0 8976 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_953
timestamp 1626908933
transform 1 0 8976 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_79
timestamp 1626908933
transform 1 0 9216 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_447
timestamp 1626908933
transform 1 0 9216 0 1 14652
box -38 -49 230 715
use L1M1_PR  L1M1_PR_163
timestamp 1626908933
transform 1 0 9456 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_951
timestamp 1626908933
transform 1 0 9456 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_463
timestamp 1626908933
transform 1 0 9504 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1032
timestamp 1626908933
transform 1 0 9504 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_113
timestamp 1626908933
transform 1 0 9408 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_743
timestamp 1626908933
transform 1 0 9408 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_46
timestamp 1626908933
transform 1 0 7584 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_21
timestamp 1626908933
transform 1 0 7584 0 1 14652
box -38 -49 1670 715
use L1M1_PR  L1M1_PR_718
timestamp 1626908933
transform 1 0 10032 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1506
timestamp 1626908933
transform 1 0 10032 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_76
timestamp 1626908933
transform 1 0 9984 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_335
timestamp 1626908933
transform 1 0 9984 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_332
timestamp 1626908933
transform 1 0 10080 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_700
timestamp 1626908933
transform 1 0 10080 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_112
timestamp 1626908933
transform 1 0 9888 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_742
timestamp 1626908933
transform 1 0 9888 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1452
timestamp 1626908933
transform 1 0 10320 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_684
timestamp 1626908933
transform 1 0 10320 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1449
timestamp 1626908933
transform 1 0 10512 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_681
timestamp 1626908933
transform 1 0 10512 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1503
timestamp 1626908933
transform 1 0 10512 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_715
timestamp 1626908933
transform 1 0 10512 0 1 14319
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_499
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_229
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_499
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_229
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_499
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_229
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_244
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_532
timestamp 1626908933
transform 1 0 10600 0 1 14652
box -200 -142 200 178
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_51
timestamp 1626908933
transform 1 0 10272 0 1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_131
timestamp 1626908933
transform 1 0 10272 0 1 14652
box -38 -49 902 715
use L1M1_PR  L1M1_PR_159
timestamp 1626908933
transform 1 0 10896 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_947
timestamp 1626908933
transform 1 0 10896 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_694
timestamp 1626908933
transform 1 0 10992 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1462
timestamp 1626908933
transform 1 0 10992 0 1 14245
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_422
timestamp 1626908933
transform 1 0 11424 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_991
timestamp 1626908933
transform 1 0 11424 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_78
timestamp 1626908933
transform 1 0 11136 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_446
timestamp 1626908933
transform 1 0 11136 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_111
timestamp 1626908933
transform 1 0 11328 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_741
timestamp 1626908933
transform 1 0 11328 0 1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_724
timestamp 1626908933
transform 1 0 11568 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1512
timestamp 1626908933
transform 1 0 11568 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_113
timestamp 1626908933
transform 1 0 11808 0 1 14652
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_33
timestamp 1626908933
transform 1 0 11808 0 1 14652
box -38 -49 902 715
use L1M1_PR  L1M1_PR_945
timestamp 1626908933
transform 1 0 11952 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_157
timestamp 1626908933
transform 1 0 11952 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1459
timestamp 1626908933
transform 1 0 11856 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_691
timestamp 1626908933
transform 1 0 11856 0 1 14245
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_740
timestamp 1626908933
transform 1 0 12672 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_110
timestamp 1626908933
transform 1 0 12672 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_962
timestamp 1626908933
transform 1 0 12768 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_393
timestamp 1626908933
transform 1 0 12768 0 1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1169
timestamp 1626908933
transform 1 0 13680 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_381
timestamp 1626908933
transform 1 0 13680 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1077
timestamp 1626908933
transform 1 0 13680 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_309
timestamp 1626908933
transform 1 0 13680 0 1 14319
box -32 -32 32 32
use osc_core_VIA3  osc_core_VIA3_7
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_2
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_7
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_2
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -28 96 28
use osc_core_VIA1  osc_core_VIA1_7
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_2
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_7
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_2
timestamp 1626908933
transform 1 0 14116 0 1 14470
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_6
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_1
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_6
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_1
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -33 96 33
use L1M1_PR  L1M1_PR_795
timestamp 1626908933
transform 1 0 14640 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_7
timestamp 1626908933
transform 1 0 14640 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_780
timestamp 1626908933
transform 1 0 14640 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_12
timestamp 1626908933
transform 1 0 14640 0 1 14319
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_228
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_516
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_484
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_214
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_484
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_214
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_484
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_214
timestamp 1626908933
transform 1 0 14600 0 1 14652
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_75
timestamp 1626908933
transform 1 0 14976 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_334
timestamp 1626908933
transform 1 0 14976 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_333
timestamp 1626908933
transform 1 0 14784 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_701
timestamp 1626908933
transform 1 0 14784 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_109
timestamp 1626908933
transform 1 0 15072 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_739
timestamp 1626908933
transform 1 0 15072 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_348
timestamp 1626908933
transform 1 0 15168 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_917
timestamp 1626908933
transform 1 0 15168 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_31
timestamp 1626908933
transform 1 0 13152 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_6
timestamp 1626908933
transform 1 0 13152 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_955
timestamp 1626908933
transform 1 0 15552 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_385
timestamp 1626908933
transform 1 0 15552 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_892
timestamp 1626908933
transform 1 0 16320 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_323
timestamp 1626908933
transform 1 0 16320 0 1 14652
box -38 -49 422 715
use M1M2_PR  M1M2_PR_45
timestamp 1626908933
transform 1 0 18000 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_813
timestamp 1626908933
transform 1 0 18000 0 1 14245
box -32 -32 32 32
use M2M3_PR  M2M3_PR_2
timestamp 1626908933
transform 1 0 18000 0 1 14189
box -33 -37 33 37
use M2M3_PR  M2M3_PR_61
timestamp 1626908933
transform 1 0 18000 0 1 14189
box -33 -37 33 37
use M3M4_PR  M3M4_PR_2
timestamp 1626908933
transform 1 0 17952 0 1 14189
box -38 -33 38 33
use M3M4_PR  M3M4_PR_23
timestamp 1626908933
transform 1 0 17952 0 1 14189
box -38 -33 38 33
use M1M2_PR  M1M2_PR_44
timestamp 1626908933
transform 1 0 18000 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_812
timestamp 1626908933
transform 1 0 18000 0 1 14837
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_359
timestamp 1626908933
transform 1 0 16704 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_929
timestamp 1626908933
transform 1 0 16704 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_41
timestamp 1626908933
transform 1 0 17472 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_16
timestamp 1626908933
transform 1 0 17472 0 1 14652
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_546
timestamp 1626908933
transform 1 0 18288 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1314
timestamp 1626908933
transform 1 0 18288 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_621
timestamp 1626908933
transform 1 0 18288 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1409
timestamp 1626908933
transform 1 0 18288 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_50
timestamp 1626908933
transform 1 0 18000 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_838
timestamp 1626908933
transform 1 0 18000 0 1 14245
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_212
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_500
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_199
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_469
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_199
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_469
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_199
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_469
timestamp 1626908933
transform 1 0 18600 0 1 14652
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_882
timestamp 1626908933
transform 1 0 19200 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_312
timestamp 1626908933
transform 1 0 19200 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_738
timestamp 1626908933
transform 1 0 19104 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_108
timestamp 1626908933
transform 1 0 19104 0 1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_904
timestamp 1626908933
transform 1 0 18960 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_116
timestamp 1626908933
transform 1 0 18960 0 1 14319
box -29 -23 29 23
use M1M2_PR  M1M2_PR_867
timestamp 1626908933
transform 1 0 19152 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_99
timestamp 1626908933
transform 1 0 19152 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_868
timestamp 1626908933
transform 1 0 20064 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_298
timestamp 1626908933
transform 1 0 20064 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_333
timestamp 1626908933
transform 1 0 19968 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_74
timestamp 1626908933
transform 1 0 19968 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_250
timestamp 1626908933
transform 1 0 21120 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_819
timestamp 1626908933
transform 1 0 21120 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_77
timestamp 1626908933
transform 1 0 20832 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_445
timestamp 1626908933
transform 1 0 20832 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_107
timestamp 1626908933
transform 1 0 21024 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_737
timestamp 1626908933
transform 1 0 21024 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_552
timestamp 1626908933
transform 1 0 21936 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1320
timestamp 1626908933
transform 1 0 21936 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_628
timestamp 1626908933
transform 1 0 21936 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1416
timestamp 1626908933
transform 1 0 21936 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_788
timestamp 1626908933
transform 1 0 22416 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_0
timestamp 1626908933
transform 1 0 22416 0 1 14097
box -29 -23 29 23
use M1M2_PR  M1M2_PR_769
timestamp 1626908933
transform 1 0 22320 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1
timestamp 1626908933
transform 1 0 22320 0 1 14097
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_454
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_184
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_454
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_184
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_454
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_184
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_484
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_196
timestamp 1626908933
transform 1 0 22600 0 1 14652
box -200 -142 200 178
use M1M2_PR  M1M2_PR_38
timestamp 1626908933
transform 1 0 22992 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_806
timestamp 1626908933
transform 1 0 22992 0 1 14319
box -32 -32 32 32
use L1M1_PR  L1M1_PR_41
timestamp 1626908933
transform 1 0 22992 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_542
timestamp 1626908933
transform 1 0 23280 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_829
timestamp 1626908933
transform 1 0 22992 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1330
timestamp 1626908933
transform 1 0 23280 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_254
timestamp 1626908933
transform 1 0 23136 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_622
timestamp 1626908933
transform 1 0 23136 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_26
timestamp 1626908933
transform 1 0 23328 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_66
timestamp 1626908933
transform 1 0 23328 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_36
timestamp 1626908933
transform 1 0 21504 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_11
timestamp 1626908933
transform 1 0 21504 0 1 14652
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_1253
timestamp 1626908933
transform 1 0 23760 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_485
timestamp 1626908933
transform 1 0 23760 0 1 14763
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1326
timestamp 1626908933
transform 1 0 23856 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_538
timestamp 1626908933
transform 1 0 23856 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1341
timestamp 1626908933
transform 1 0 24048 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_553
timestamp 1626908933
transform 1 0 24048 0 1 14763
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_332
timestamp 1626908933
transform 1 0 24096 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_73
timestamp 1626908933
transform 1 0 24096 0 1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1294
timestamp 1626908933
transform 1 0 24048 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_506
timestamp 1626908933
transform 1 0 24048 0 1 14245
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1215
timestamp 1626908933
transform 1 0 24144 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_447
timestamp 1626908933
transform 1 0 24144 0 1 14245
box -32 -32 32 32
use L1M1_PR  L1M1_PR_504
timestamp 1626908933
transform 1 0 24240 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1292
timestamp 1626908933
transform 1 0 24240 0 1 14245
box -29 -23 29 23
use L1M1_PR  L1M1_PR_479
timestamp 1626908933
transform 1 0 24624 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1267
timestamp 1626908933
transform 1 0 24624 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__nand3_4  sky130_fd_sc_hs__nand3_4_1
timestamp 1626908933
transform 1 0 24192 0 1 14652
box -38 -49 1286 715
use sky130_fd_sc_hs__nand3_4  sky130_fd_sc_hs__nand3_4_3
timestamp 1626908933
transform 1 0 24192 0 1 14652
box -38 -49 1286 715
use M1M2_PR  M1M2_PR_405
timestamp 1626908933
transform 1 0 24912 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1173
timestamp 1626908933
transform 1 0 24912 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_440
timestamp 1626908933
transform 1 0 25488 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_469
timestamp 1626908933
transform 1 0 25776 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1208
timestamp 1626908933
transform 1 0 25488 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1237
timestamp 1626908933
transform 1 0 25776 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_446
timestamp 1626908933
transform 1 0 24912 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1214
timestamp 1626908933
transform 1 0 24912 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_442
timestamp 1626908933
transform 1 0 25680 0 1 14541
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1210
timestamp 1626908933
transform 1 0 25680 0 1 14541
box -32 -32 32 32
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_31
timestamp 1626908933
transform 1 0 25440 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__dlygate4sd3_1  sky130_fd_sc_hs__dlygate4sd3_1_71
timestamp 1626908933
transform 1 0 25440 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_702
timestamp 1626908933
transform 1 0 26208 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_334
timestamp 1626908933
transform 1 0 26208 0 1 14652
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1222
timestamp 1626908933
transform 1 0 26928 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_434
timestamp 1626908933
transform 1 0 26928 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1225
timestamp 1626908933
transform 1 0 26736 0 1 14393
box -29 -23 29 23
use L1M1_PR  L1M1_PR_437
timestamp 1626908933
transform 1 0 26736 0 1 14393
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1130
timestamp 1626908933
transform 1 0 26640 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_362
timestamp 1626908933
transform 1 0 26640 0 1 14319
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_169
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_439
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_169
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_439
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_169
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_439
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -49 200 49
use L1M1_PR  L1M1_PR_442
timestamp 1626908933
transform 1 0 26928 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1230
timestamp 1626908933
transform 1 0 26928 0 1 14763
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_468
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_180
timestamp 1626908933
transform 1 0 26600 0 1 14652
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1190
timestamp 1626908933
transform 1 0 26400 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_560
timestamp 1626908933
transform 1 0 26400 0 1 14652
box -38 -49 134 715
use M1M2_PR  M1M2_PR_473
timestamp 1626908933
transform 1 0 27024 0 1 14171
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1241
timestamp 1626908933
transform 1 0 27024 0 1 14171
box -32 -32 32 32
use L1M1_PR  L1M1_PR_436
timestamp 1626908933
transform 1 0 27024 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1224
timestamp 1626908933
transform 1 0 27024 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_501
timestamp 1626908933
transform 1 0 27216 0 1 14541
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1289
timestamp 1626908933
transform 1 0 27216 0 1 14541
box -29 -23 29 23
use M1M2_PR  M1M2_PR_372
timestamp 1626908933
transform 1 0 27216 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1140
timestamp 1626908933
transform 1 0 27216 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_377
timestamp 1626908933
transform 1 0 27120 0 1 14837
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1145
timestamp 1626908933
transform 1 0 27120 0 1 14837
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_703
timestamp 1626908933
transform 1 0 27264 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_335
timestamp 1626908933
transform 1 0 27264 0 1 14652
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1143
timestamp 1626908933
transform 1 0 27408 0 1 14245
box -32 -32 32 32
use M1M2_PR  M1M2_PR_375
timestamp 1626908933
transform 1 0 27408 0 1 14245
box -32 -32 32 32
use sky130_fd_sc_hs__and4_2  sky130_fd_sc_hs__and4_2_1
timestamp 1626908933
transform -1 0 27264 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__and4_2  sky130_fd_sc_hs__and4_2_4
timestamp 1626908933
transform -1 0 27264 0 1 14652
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1193
timestamp 1626908933
transform 1 0 29040 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_425
timestamp 1626908933
transform 1 0 29040 0 1 14319
box -32 -32 32 32
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_23
timestamp 1626908933
transform 1 0 27456 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_7
timestamp 1626908933
transform 1 0 27456 0 1 14652
box -38 -49 1670 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_76
timestamp 1626908933
transform 1 0 29088 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_444
timestamp 1626908933
transform 1 0 29088 0 1 14652
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1271
timestamp 1626908933
transform 1 0 29808 0 1 14097
box -29 -23 29 23
use L1M1_PR  L1M1_PR_483
timestamp 1626908933
transform 1 0 29808 0 1 14097
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1177
timestamp 1626908933
transform 1 0 29904 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_409
timestamp 1626908933
transform 1 0 29904 0 1 14319
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1178
timestamp 1626908933
transform 1 0 29712 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_410
timestamp 1626908933
transform 1 0 29712 0 1 14097
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1176
timestamp 1626908933
transform 1 0 29904 0 1 14763
box -32 -32 32 32
use M1M2_PR  M1M2_PR_408
timestamp 1626908933
transform 1 0 29904 0 1 14763
box -32 -32 32 32
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_5
timestamp 1626908933
transform 1 0 29664 0 1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_0
timestamp 1626908933
transform 1 0 29664 0 1 14652
box -38 -49 326 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_128
timestamp 1626908933
transform 1 0 29280 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_697
timestamp 1626908933
transform 1 0 29280 0 1 14652
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1269
timestamp 1626908933
transform 1 0 29904 0 1 14763
box -29 -23 29 23
use L1M1_PR  L1M1_PR_481
timestamp 1626908933
transform 1 0 29904 0 1 14763
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_331
timestamp 1626908933
transform 1 0 29952 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_72
timestamp 1626908933
transform 1 0 29952 0 1 14652
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1270
timestamp 1626908933
transform 1 0 29904 0 1 14319
box -29 -23 29 23
use L1M1_PR  L1M1_PR_482
timestamp 1626908933
transform 1 0 29904 0 1 14319
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_736
timestamp 1626908933
transform 1 0 30240 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_106
timestamp 1626908933
transform 1 0 30240 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_443
timestamp 1626908933
transform 1 0 30048 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_75
timestamp 1626908933
transform 1 0 30048 0 1 14652
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_154
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_424
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_154
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_424
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_154
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_424
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_164
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_452
timestamp 1626908933
transform 1 0 30600 0 1 14652
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_112
timestamp 1626908933
transform 1 0 30336 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_682
timestamp 1626908933
transform 1 0 30336 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_442
timestamp 1626908933
transform 1 0 31104 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_74
timestamp 1626908933
transform 1 0 31104 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_660
timestamp 1626908933
transform 1 0 31296 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_91
timestamp 1626908933
transform 1 0 31296 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_652
timestamp 1626908933
transform 1 0 31680 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_82
timestamp 1626908933
transform 1 0 31680 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_735
timestamp 1626908933
transform 1 0 32448 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_105
timestamp 1626908933
transform 1 0 32448 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_627
timestamp 1626908933
transform 1 0 32544 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_58
timestamp 1626908933
transform 1 0 32544 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_622
timestamp 1626908933
transform 1 0 32928 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_52
timestamp 1626908933
transform 1 0 32928 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_734
timestamp 1626908933
transform 1 0 33696 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_104
timestamp 1626908933
transform 1 0 33696 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_594
timestamp 1626908933
transform 1 0 33792 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_25
timestamp 1626908933
transform 1 0 33792 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_592
timestamp 1626908933
transform 1 0 34176 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_22
timestamp 1626908933
transform 1 0 34176 0 1 14652
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_409
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_139
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_409
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_139
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_409
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_139
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_148
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_436
timestamp 1626908933
transform 1 0 34600 0 1 14652
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_71
timestamp 1626908933
transform 1 0 34944 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_330
timestamp 1626908933
transform 1 0 34944 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_4
timestamp 1626908933
transform 1 0 35040 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_573
timestamp 1626908933
transform 1 0 35040 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_336
timestamp 1626908933
transform 1 0 35424 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_704
timestamp 1626908933
transform 1 0 35424 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_561
timestamp 1626908933
transform 1 0 35616 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1191
timestamp 1626908933
transform 1 0 35616 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_441
timestamp 1626908933
transform 1 0 288 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_73
timestamp 1626908933
transform 1 0 288 0 -1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_291
timestamp 1626908933
transform 1 0 624 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1059
timestamp 1626908933
transform 1 0 624 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_355
timestamp 1626908933
transform 1 0 816 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1143
timestamp 1626908933
transform 1 0 816 0 1 14985
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_420
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_132
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_123
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_393
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_123
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_393
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_123
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_393
timestamp 1626908933
transform 1 0 600 0 1 15318
box -200 -49 200 49
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_95
timestamp 1626908933
transform -1 0 1344 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_40
timestamp 1626908933
transform -1 0 1344 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_567
timestamp 1626908933
transform 1 0 480 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1136
timestamp 1626908933
transform 1 0 480 0 -1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_154
timestamp 1626908933
transform 1 0 1008 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_922
timestamp 1626908933
transform 1 0 1008 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_197
timestamp 1626908933
transform 1 0 1008 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_985
timestamp 1626908933
transform 1 0 1008 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_153
timestamp 1626908933
transform 1 0 1008 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_921
timestamp 1626908933
transform 1 0 1008 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_293
timestamp 1626908933
transform 1 0 1296 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1061
timestamp 1626908933
transform 1 0 1296 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_360
timestamp 1626908933
transform 1 0 1296 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1148
timestamp 1626908933
transform 1 0 1296 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_337
timestamp 1626908933
transform 1 0 1344 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_705
timestamp 1626908933
transform 1 0 1344 0 -1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_191
timestamp 1626908933
transform 1 0 1488 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_979
timestamp 1626908933
transform 1 0 1488 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_98
timestamp 1626908933
transform 1 0 1536 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_43
timestamp 1626908933
transform 1 0 1536 0 -1 15984
box -38 -49 518 715
use L1M1_PR  L1M1_PR_976
timestamp 1626908933
transform 1 0 1968 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_188
timestamp 1626908933
transform 1 0 1968 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1141
timestamp 1626908933
transform 1 0 2064 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_353
timestamp 1626908933
transform 1 0 2064 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1417
timestamp 1626908933
transform 1 0 2160 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_649
timestamp 1626908933
transform 1 0 2160 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1056
timestamp 1626908933
transform 1 0 2064 0 1 15133
box -32 -32 32 32
use M1M2_PR  M1M2_PR_288
timestamp 1626908933
transform 1 0 2064 0 1 15133
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_329
timestamp 1626908933
transform 1 0 2496 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_70
timestamp 1626908933
transform 1 0 2496 0 -1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1152
timestamp 1626908933
transform 1 0 2256 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_384
timestamp 1626908933
transform 1 0 2256 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1467
timestamp 1626908933
transform 1 0 2352 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1238
timestamp 1626908933
transform 1 0 2448 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_679
timestamp 1626908933
transform 1 0 2352 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_450
timestamp 1626908933
transform 1 0 2448 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_36
timestamp 1626908933
transform 1 0 2016 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_91
timestamp 1626908933
transform 1 0 2016 0 -1 15984
box -38 -49 518 715
use L1M1_PR  L1M1_PR_344
timestamp 1626908933
transform 1 0 2544 0 1 14837
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1132
timestamp 1626908933
transform 1 0 2544 0 1 14837
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_538
timestamp 1626908933
transform 1 0 2688 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1107
timestamp 1626908933
transform 1 0 2688 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_103
timestamp 1626908933
transform 1 0 2592 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_733
timestamp 1626908933
transform 1 0 2592 0 -1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_319
timestamp 1626908933
transform 1 0 3504 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1087
timestamp 1626908933
transform 1 0 3504 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_392
timestamp 1626908933
transform 1 0 3504 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1180
timestamp 1626908933
transform 1 0 3504 0 1 14985
box -29 -23 29 23
use M3M4_PR  M3M4_PR_15
timestamp 1626908933
transform 1 0 3552 0 1 15043
box -38 -33 38 33
use M3M4_PR  M3M4_PR_36
timestamp 1626908933
transform 1 0 3552 0 1 15043
box -38 -33 38 33
use M2M3_PR  M2M3_PR_15
timestamp 1626908933
transform 1 0 3696 0 1 15043
box -33 -37 33 37
use M2M3_PR  M2M3_PR_74
timestamp 1626908933
transform 1 0 3696 0 1 15043
box -33 -37 33 37
use M1M2_PR  M1M2_PR_568
timestamp 1626908933
transform 1 0 3312 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1336
timestamp 1626908933
transform 1 0 3312 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_144
timestamp 1626908933
transform 1 0 3696 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_912
timestamp 1626908933
transform 1 0 3696 0 1 15059
box -32 -32 32 32
use L1M1_PR  L1M1_PR_181
timestamp 1626908933
transform 1 0 3696 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_969
timestamp 1626908933
transform 1 0 3696 0 1 15059
box -29 -23 29 23
use M1M2_PR  M1M2_PR_146
timestamp 1626908933
transform 1 0 3600 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_914
timestamp 1626908933
transform 1 0 3600 0 1 15577
box -32 -32 32 32
use L1M1_PR  L1M1_PR_183
timestamp 1626908933
transform 1 0 3600 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_971
timestamp 1626908933
transform 1 0 3600 0 1 15577
box -29 -23 29 23
use M2M3_PR  M2M3_PR_17
timestamp 1626908933
transform 1 0 3600 0 1 15531
box -33 -37 33 37
use M2M3_PR  M2M3_PR_76
timestamp 1626908933
transform 1 0 3600 0 1 15531
box -33 -37 33 37
use M3M4_PR  M3M4_PR_14
timestamp 1626908933
transform 1 0 3552 0 1 15531
box -38 -33 38 33
use M3M4_PR  M3M4_PR_35
timestamp 1626908933
transform 1 0 3552 0 1 15531
box -38 -33 38 33
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_25
timestamp 1626908933
transform 1 0 3072 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_0
timestamp 1626908933
transform 1 0 3072 0 -1 15984
box -38 -49 1670 715
use L1M1_PR  L1M1_PR_892
timestamp 1626908933
transform 1 0 4560 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_104
timestamp 1626908933
transform 1 0 4560 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_857
timestamp 1626908933
transform 1 0 4560 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_89
timestamp 1626908933
transform 1 0 4560 0 1 14985
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_378
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_108
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_378
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_108
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_378
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_108
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_404
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_116
timestamp 1626908933
transform 1 0 4600 0 1 15318
box -200 -142 200 178
use L1M1_PR  L1M1_PR_961
timestamp 1626908933
transform 1 0 4560 0 1 15503
box -29 -23 29 23
use L1M1_PR  L1M1_PR_173
timestamp 1626908933
transform 1 0 4560 0 1 15503
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_562
timestamp 1626908933
transform 1 0 4704 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1192
timestamp 1626908933
transform 1 0 4704 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_47
timestamp 1626908933
transform 1 0 4800 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_127
timestamp 1626908933
transform 1 0 4800 0 -1 15984
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1128
timestamp 1626908933
transform 1 0 5232 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_340
timestamp 1626908933
transform 1 0 5232 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1048
timestamp 1626908933
transform 1 0 5136 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_280
timestamp 1626908933
transform 1 0 5136 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_883
timestamp 1626908933
transform 1 0 5424 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_95
timestamp 1626908933
transform 1 0 5424 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1558
timestamp 1626908933
transform 1 0 6000 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_770
timestamp 1626908933
transform 1 0 6000 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1509
timestamp 1626908933
transform 1 0 6000 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_741
timestamp 1626908933
transform 1 0 6000 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_62
timestamp 1626908933
transform 1 0 5664 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_142
timestamp 1626908933
transform 1 0 5664 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_139
timestamp 1626908933
transform 1 0 6528 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_59
timestamp 1626908933
transform 1 0 6528 0 -1 15984
box -38 -49 902 715
use L1M1_PR  L1M1_PR_820
timestamp 1626908933
transform 1 0 6384 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_32
timestamp 1626908933
transform 1 0 6384 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_798
timestamp 1626908933
transform 1 0 6288 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_30
timestamp 1626908933
transform 1 0 6288 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_563
timestamp 1626908933
transform 1 0 7392 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1193
timestamp 1626908933
transform 1 0 7392 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_69
timestamp 1626908933
transform 1 0 7488 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_328
timestamp 1626908933
transform 1 0 7488 0 -1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_110
timestamp 1626908933
transform 1 0 8112 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_878
timestamp 1626908933
transform 1 0 8112 0 1 15059
box -32 -32 32 32
use L1M1_PR  L1M1_PR_129
timestamp 1626908933
transform 1 0 8112 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_917
timestamp 1626908933
transform 1 0 8112 0 1 15059
box -29 -23 29 23
use M2M3_PR  M2M3_PR_8
timestamp 1626908933
transform 1 0 8112 0 1 15043
box -33 -37 33 37
use M2M3_PR  M2M3_PR_67
timestamp 1626908933
transform 1 0 8112 0 1 15043
box -33 -37 33 37
use M3M4_PR  M3M4_PR_7
timestamp 1626908933
transform 1 0 8112 0 1 15043
box -38 -33 38 33
use M3M4_PR  M3M4_PR_28
timestamp 1626908933
transform 1 0 8112 0 1 15043
box -38 -33 38 33
use M1M2_PR  M1M2_PR_314
timestamp 1626908933
transform 1 0 8304 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1082
timestamp 1626908933
transform 1 0 8304 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_386
timestamp 1626908933
transform 1 0 8304 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1174
timestamp 1626908933
transform 1 0 8304 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_952
timestamp 1626908933
transform 1 0 8976 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_164
timestamp 1626908933
transform 1 0 8976 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_898
timestamp 1626908933
transform 1 0 8976 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_130
timestamp 1626908933
transform 1 0 8976 0 1 14985
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_363
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_93
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_363
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_93
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_363
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_93
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_388
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_100
timestamp 1626908933
transform 1 0 8600 0 1 15318
box -200 -142 200 178
use M1M2_PR  M1M2_PR_566
timestamp 1626908933
transform 1 0 9648 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1334
timestamp 1626908933
transform 1 0 9648 0 1 15207
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_564
timestamp 1626908933
transform 1 0 9216 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1194
timestamp 1626908933
transform 1 0 9216 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_126
timestamp 1626908933
transform 1 0 9072 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_914
timestamp 1626908933
transform 1 0 9072 0 1 15429
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_57
timestamp 1626908933
transform 1 0 9312 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_137
timestamp 1626908933
transform 1 0 9312 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_45
timestamp 1626908933
transform 1 0 7584 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_20
timestamp 1626908933
transform 1 0 7584 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_338
timestamp 1626908933
transform 1 0 10176 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_706
timestamp 1626908933
transform 1 0 10176 0 -1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_577
timestamp 1626908933
transform 1 0 10320 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_683
timestamp 1626908933
transform 1 0 10320 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1345
timestamp 1626908933
transform 1 0 10320 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1451
timestamp 1626908933
transform 1 0 10320 0 1 15059
box -32 -32 32 32
use L1M1_PR  L1M1_PR_714
timestamp 1626908933
transform 1 0 10512 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1502
timestamp 1626908933
transform 1 0 10512 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_58
timestamp 1626908933
transform 1 0 10368 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_138
timestamp 1626908933
transform 1 0 10368 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_116
timestamp 1626908933
transform 1 0 11520 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_36
timestamp 1626908933
transform 1 0 11520 0 -1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1195
timestamp 1626908933
transform 1 0 11424 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_565
timestamp 1626908933
transform 1 0 11424 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_707
timestamp 1626908933
transform 1 0 11232 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_339
timestamp 1626908933
transform 1 0 11232 0 -1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_948
timestamp 1626908933
transform 1 0 10800 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_160
timestamp 1626908933
transform 1 0 10800 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_709
timestamp 1626908933
transform 1 0 11952 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1497
timestamp 1626908933
transform 1 0 11952 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_70
timestamp 1626908933
transform 1 0 12240 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_838
timestamp 1626908933
transform 1 0 12240 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_566
timestamp 1626908933
transform 1 0 12384 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1196
timestamp 1626908933
transform 1 0 12384 0 -1 15984
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_372
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_84
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_78
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_348
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_78
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_348
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_78
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_348
timestamp 1626908933
transform 1 0 12600 0 1 15318
box -200 -49 200 49
use L1M1_PR  L1M1_PR_80
timestamp 1626908933
transform 1 0 12528 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_868
timestamp 1626908933
transform 1 0 12528 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_392
timestamp 1626908933
transform 1 0 12768 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_961
timestamp 1626908933
transform 1 0 12768 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_72
timestamp 1626908933
transform 1 0 12576 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_440
timestamp 1626908933
transform 1 0 12576 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_68
timestamp 1626908933
transform 1 0 12480 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_327
timestamp 1626908933
transform 1 0 12480 0 -1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_67
timestamp 1626908933
transform 1 0 13104 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_835
timestamp 1626908933
transform 1 0 13104 0 1 14985
box -32 -32 32 32
use M2M3_PR  M2M3_PR_4
timestamp 1626908933
transform 1 0 13104 0 1 15043
box -33 -37 33 37
use M2M3_PR  M2M3_PR_63
timestamp 1626908933
transform 1 0 13104 0 1 15043
box -33 -37 33 37
use M1M2_PR  M1M2_PR_308
timestamp 1626908933
transform 1 0 13680 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1076
timestamp 1626908933
transform 1 0 13680 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_380
timestamp 1626908933
transform 1 0 13680 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1168
timestamp 1626908933
transform 1 0 13680 0 1 14985
box -29 -23 29 23
use M3M4_PR  M3M4_PR_5
timestamp 1626908933
transform 1 0 14112 0 1 15043
box -38 -33 38 33
use M3M4_PR  M3M4_PR_26
timestamp 1626908933
transform 1 0 14112 0 1 15043
box -38 -33 38 33
use osc_core_VIA2  osc_core_VIA2_1
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_6
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_1
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_6
timestamp 1626908933
transform 1 0 14116 0 1 14834
box -97 -28 96 28
use M1M2_PR  M1M2_PR_17
timestamp 1626908933
transform 1 0 14544 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_785
timestamp 1626908933
transform 1 0 14544 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_10
timestamp 1626908933
transform 1 0 14928 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_778
timestamp 1626908933
transform 1 0 14928 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_11
timestamp 1626908933
transform 1 0 14544 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_799
timestamp 1626908933
transform 1 0 14544 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_71
timestamp 1626908933
transform 1 0 14784 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_439
timestamp 1626908933
transform 1 0 14784 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_406
timestamp 1626908933
transform 1 0 14976 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_976
timestamp 1626908933
transform 1 0 14976 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_30
timestamp 1626908933
transform 1 0 13152 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_5
timestamp 1626908933
transform 1 0 13152 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_342
timestamp 1626908933
transform 1 0 15840 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_911
timestamp 1626908933
transform 1 0 15840 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_102
timestamp 1626908933
transform 1 0 15744 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_732
timestamp 1626908933
transform 1 0 15744 0 -1 15984
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_68
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_356
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_63
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_333
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_63
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_333
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_63
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_333
timestamp 1626908933
transform 1 0 16600 0 1 15318
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_377
timestamp 1626908933
transform 1 0 16224 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_947
timestamp 1626908933
transform 1 0 16224 0 -1 15984
box -38 -49 806 715
use M1M2_PR  M1M2_PR_575
timestamp 1626908933
transform 1 0 16848 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1343
timestamp 1626908933
transform 1 0 16848 0 1 15207
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_318
timestamp 1626908933
transform 1 0 16992 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_887
timestamp 1626908933
transform 1 0 16992 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_67
timestamp 1626908933
transform 1 0 17376 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_326
timestamp 1626908933
transform 1 0 17376 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_624
timestamp 1626908933
transform 1 0 17904 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1412
timestamp 1626908933
transform 1 0 17904 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_105
timestamp 1626908933
transform 1 0 17808 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_873
timestamp 1626908933
transform 1 0 17808 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_43
timestamp 1626908933
transform 1 0 18000 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_811
timestamp 1626908933
transform 1 0 18000 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_40
timestamp 1626908933
transform 1 0 17472 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_15
timestamp 1626908933
transform 1 0 17472 0 -1 15984
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_545
timestamp 1626908933
transform 1 0 18288 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1313
timestamp 1626908933
transform 1 0 18288 0 1 14911
box -32 -32 32 32
use L1M1_PR  L1M1_PR_47
timestamp 1626908933
transform 1 0 18384 0 1 14837
box -29 -23 29 23
use L1M1_PR  L1M1_PR_835
timestamp 1626908933
transform 1 0 18384 0 1 14837
box -29 -23 29 23
use M1M2_PR  M1M2_PR_103
timestamp 1626908933
transform 1 0 18672 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_871
timestamp 1626908933
transform 1 0 18672 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_49
timestamp 1626908933
transform 1 0 18000 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_837
timestamp 1626908933
transform 1 0 18000 0 1 15577
box -29 -23 29 23
use M1M2_PR  M1M2_PR_102
timestamp 1626908933
transform 1 0 18672 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_870
timestamp 1626908933
transform 1 0 18672 0 1 15503
box -32 -32 32 32
use M1M2_PR  M1M2_PR_98
timestamp 1626908933
transform 1 0 19152 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_866
timestamp 1626908933
transform 1 0 19152 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_115
timestamp 1626908933
transform 1 0 18960 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_903
timestamp 1626908933
transform 1 0 18960 0 1 14985
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_70
timestamp 1626908933
transform 1 0 19104 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_438
timestamp 1626908933
transform 1 0 19104 0 -1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_46
timestamp 1626908933
transform 1 0 18960 0 1 15503
box -29 -23 29 23
use L1M1_PR  L1M1_PR_834
timestamp 1626908933
transform 1 0 18960 0 1 15503
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_101
timestamp 1626908933
transform 1 0 19296 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_731
timestamp 1626908933
transform 1 0 19296 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_311
timestamp 1626908933
transform 1 0 19392 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_881
timestamp 1626908933
transform 1 0 19392 0 -1 15984
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_340
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_52
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_318
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_48
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_318
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_48
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_318
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_48
timestamp 1626908933
transform 1 0 20600 0 1 15318
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_730
timestamp 1626908933
transform 1 0 20160 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_100
timestamp 1626908933
transform 1 0 20160 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_265
timestamp 1626908933
transform 1 0 20256 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_834
timestamp 1626908933
transform 1 0 20256 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_856
timestamp 1626908933
transform 1 0 20640 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_286
timestamp 1626908933
transform 1 0 20640 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_325
timestamp 1626908933
transform 1 0 21408 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_66
timestamp 1626908933
transform 1 0 21408 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1415
timestamp 1626908933
transform 1 0 21936 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_627
timestamp 1626908933
transform 1 0 21936 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1319
timestamp 1626908933
transform 1 0 21936 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_551
timestamp 1626908933
transform 1 0 21936 0 1 14985
box -32 -32 32 32
use M3M4_PR  M3M4_PR_21
timestamp 1626908933
transform 1 0 22224 0 1 15043
box -38 -33 38 33
use M3M4_PR  M3M4_PR_0
timestamp 1626908933
transform 1 0 22224 0 1 15043
box -38 -33 38 33
use M2M3_PR  M2M3_PR_60
timestamp 1626908933
transform 1 0 22224 0 1 15043
box -33 -37 33 37
use M2M3_PR  M2M3_PR_1
timestamp 1626908933
transform 1 0 22224 0 1 15043
box -33 -37 33 37
use L1M1_PR  L1M1_PR_792
timestamp 1626908933
transform 1 0 22224 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_4
timestamp 1626908933
transform 1 0 22224 0 1 15059
box -29 -23 29 23
use M1M2_PR  M1M2_PR_772
timestamp 1626908933
transform 1 0 22224 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_4
timestamp 1626908933
transform 1 0 22224 0 1 15059
box -32 -32 32 32
use L1M1_PR  L1M1_PR_791
timestamp 1626908933
transform 1 0 22224 0 1 15577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3
timestamp 1626908933
transform 1 0 22224 0 1 15577
box -29 -23 29 23
use M1M2_PR  M1M2_PR_771
timestamp 1626908933
transform 1 0 22224 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3
timestamp 1626908933
transform 1 0 22224 0 1 15577
box -32 -32 32 32
use L1M1_PR  L1M1_PR_828
timestamp 1626908933
transform 1 0 22992 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_40
timestamp 1626908933
transform 1 0 22992 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1263
timestamp 1626908933
transform 1 0 22896 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_805
timestamp 1626908933
transform 1 0 22992 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_495
timestamp 1626908933
transform 1 0 22896 0 1 15059
box -32 -32 32 32
use M1M2_PR  M1M2_PR_37
timestamp 1626908933
transform 1 0 22992 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_437
timestamp 1626908933
transform 1 0 23136 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_69
timestamp 1626908933
transform 1 0 23136 0 -1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_1259
timestamp 1626908933
transform 1 0 23280 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_491
timestamp 1626908933
transform 1 0 23280 0 1 14911
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1347
timestamp 1626908933
transform 1 0 23376 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_559
timestamp 1626908933
transform 1 0 23376 0 1 14911
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_244
timestamp 1626908933
transform 1 0 23328 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_814
timestamp 1626908933
transform 1 0 23328 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_35
timestamp 1626908933
transform 1 0 21504 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__nand2_8  sky130_fd_sc_hs__nand2_8_10
timestamp 1626908933
transform 1 0 21504 0 -1 15984
box -38 -49 1670 715
use M1M2_PR  M1M2_PR_361
timestamp 1626908933
transform 1 0 24144 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_429
timestamp 1626908933
transform 1 0 24048 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1129
timestamp 1626908933
transform 1 0 24144 0 1 15207
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1197
timestamp 1626908933
transform 1 0 24048 0 1 14985
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_567
timestamp 1626908933
transform 1 0 24096 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1197
timestamp 1626908933
transform 1 0 24096 0 -1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1281
timestamp 1626908933
transform 1 0 24432 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_493
timestamp 1626908933
transform 1 0 24432 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1175
timestamp 1626908933
transform 1 0 24720 0 1 15133
box -32 -32 32 32
use M1M2_PR  M1M2_PR_407
timestamp 1626908933
transform 1 0 24720 0 1 15133
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1291
timestamp 1626908933
transform 1 0 24816 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_503
timestamp 1626908933
transform 1 0 24816 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_432
timestamp 1626908933
transform 1 0 24336 0 1 15207
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1220
timestamp 1626908933
transform 1 0 24336 0 1 15207
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_33
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_303
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_33
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_303
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_33
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_303
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_324
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_36
timestamp 1626908933
transform 1 0 24600 0 1 15318
box -200 -142 200 178
use sky130_fd_sc_hs__nand3_4  sky130_fd_sc_hs__nand3_4_0
timestamp 1626908933
transform 1 0 24192 0 -1 15984
box -38 -49 1286 715
use sky130_fd_sc_hs__nand3_4  sky130_fd_sc_hs__nand3_4_2
timestamp 1626908933
transform 1 0 24192 0 -1 15984
box -38 -49 1286 715
use L1M1_PR  L1M1_PR_1298
timestamp 1626908933
transform 1 0 25200 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_510
timestamp 1626908933
transform 1 0 25200 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1221
timestamp 1626908933
transform 1 0 25200 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_453
timestamp 1626908933
transform 1 0 25200 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1213
timestamp 1626908933
transform 1 0 24912 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_445
timestamp 1626908933
transform 1 0 24912 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1212
timestamp 1626908933
transform 1 0 25008 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_444
timestamp 1626908933
transform 1 0 25008 0 1 15577
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_765
timestamp 1626908933
transform 1 0 25440 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_196
timestamp 1626908933
transform 1 0 25440 0 -1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_499
timestamp 1626908933
transform 1 0 25584 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1267
timestamp 1626908933
transform 1 0 25584 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_572
timestamp 1626908933
transform 1 0 25584 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1360
timestamp 1626908933
transform 1 0 25584 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_565
timestamp 1626908933
transform 1 0 26160 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1353
timestamp 1626908933
transform 1 0 26160 0 1 15059
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_200
timestamp 1626908933
transform 1 0 25824 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_770
timestamp 1626908933
transform 1 0 25824 0 -1 15984
box -38 -49 806 715
use L1M1_PR  L1M1_PR_443
timestamp 1626908933
transform 1 0 26832 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_492
timestamp 1626908933
transform 1 0 26640 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1231
timestamp 1626908933
transform 1 0 26832 0 1 14911
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1280
timestamp 1626908933
transform 1 0 26640 0 1 14911
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1144
timestamp 1626908933
transform 1 0 27120 0 1 15577
box -32 -32 32 32
use M1M2_PR  M1M2_PR_376
timestamp 1626908933
transform 1 0 27120 0 1 15577
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1233
timestamp 1626908933
transform 1 0 27024 0 1 14837
box -29 -23 29 23
use L1M1_PR  L1M1_PR_445
timestamp 1626908933
transform 1 0 27024 0 1 14837
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1232
timestamp 1626908933
transform 1 0 27312 0 1 15059
box -29 -23 29 23
use L1M1_PR  L1M1_PR_444
timestamp 1626908933
transform 1 0 27312 0 1 15059
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_324
timestamp 1626908933
transform 1 0 27360 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_65
timestamp 1626908933
transform 1 0 27360 0 -1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1142
timestamp 1626908933
transform 1 0 27408 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_374
timestamp 1626908933
transform 1 0 27408 0 1 14911
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_178
timestamp 1626908933
transform 1 0 26592 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_748
timestamp 1626908933
transform 1 0 26592 0 -1 15984
box -38 -49 806 715
use M1M2_PR  M1M2_PR_424
timestamp 1626908933
transform 1 0 29040 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1192
timestamp 1626908933
transform 1 0 29040 0 1 14911
box -32 -32 32 32
use M1M2_PR  M1M2_PR_640
timestamp 1626908933
transform 1 0 28080 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1408
timestamp 1626908933
transform 1 0 28080 0 1 15429
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_20
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_308
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_18
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_288
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_18
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_288
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_18
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_288
timestamp 1626908933
transform 1 0 28600 0 1 15318
box -200 -49 200 49
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_22
timestamp 1626908933
transform 1 0 27456 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__inv_16  sky130_fd_sc_hs__inv_16_6
timestamp 1626908933
transform 1 0 27456 0 -1 15984
box -38 -49 1670 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_340
timestamp 1626908933
transform 1 0 29472 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_708
timestamp 1626908933
transform 1 0 29472 0 -1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1266
timestamp 1626908933
transform 1 0 29808 0 1 14985
box -29 -23 29 23
use L1M1_PR  L1M1_PR_478
timestamp 1626908933
transform 1 0 29808 0 1 14985
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1172
timestamp 1626908933
transform 1 0 29808 0 1 14985
box -32 -32 32 32
use M1M2_PR  M1M2_PR_404
timestamp 1626908933
transform 1 0 29808 0 1 14985
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1460
timestamp 1626908933
transform 1 0 29616 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_672
timestamp 1626908933
transform 1 0 29616 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1265
timestamp 1626908933
transform 1 0 29808 0 1 15429
box -29 -23 29 23
use L1M1_PR  L1M1_PR_477
timestamp 1626908933
transform 1 0 29808 0 1 15429
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1171
timestamp 1626908933
transform 1 0 29808 0 1 15429
box -32 -32 32 32
use M1M2_PR  M1M2_PR_403
timestamp 1626908933
transform 1 0 29808 0 1 15429
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_26
timestamp 1626908933
transform 1 0 29664 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_6
timestamp 1626908933
transform 1 0 29664 0 -1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_6
timestamp 1626908933
transform 1 0 29088 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_15
timestamp 1626908933
transform 1 0 29088 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_436
timestamp 1626908933
transform 1 0 30144 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_68
timestamp 1626908933
transform 1 0 30144 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_681
timestamp 1626908933
transform 1 0 30336 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_111
timestamp 1626908933
transform 1 0 30336 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_435
timestamp 1626908933
transform 1 0 31104 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_67
timestamp 1626908933
transform 1 0 31104 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_659
timestamp 1626908933
transform 1 0 31296 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_90
timestamp 1626908933
transform 1 0 31296 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_651
timestamp 1626908933
transform 1 0 31680 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_81
timestamp 1626908933
transform 1 0 31680 0 -1 15984
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_292
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_4
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_273
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_3
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_273
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_3
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_273
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_3
timestamp 1626908933
transform 1 0 32600 0 1 15318
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_323
timestamp 1626908933
transform 1 0 32448 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_64
timestamp 1626908933
transform 1 0 32448 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_57
timestamp 1626908933
transform 1 0 32544 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_626
timestamp 1626908933
transform 1 0 32544 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_621
timestamp 1626908933
transform 1 0 32928 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_51
timestamp 1626908933
transform 1 0 32928 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_729
timestamp 1626908933
transform 1 0 33696 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_99
timestamp 1626908933
transform 1 0 33696 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_593
timestamp 1626908933
transform 1 0 33792 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_24
timestamp 1626908933
transform 1 0 33792 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_591
timestamp 1626908933
transform 1 0 34176 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_21
timestamp 1626908933
transform 1 0 34176 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_3
timestamp 1626908933
transform 1 0 34944 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_573
timestamp 1626908933
transform 1 0 34944 0 -1 15984
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1413
timestamp 1626908933
transform 1 0 48 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_645
timestamp 1626908933
transform 1 0 48 0 1 15873
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_322
timestamp 1626908933
transform 1 0 288 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_63
timestamp 1626908933
transform 1 0 288 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1135
timestamp 1626908933
transform 1 0 480 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_566
timestamp 1626908933
transform 1 0 480 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_727
timestamp 1626908933
transform 1 0 864 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_97
timestamp 1626908933
transform 1 0 864 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_728
timestamp 1626908933
transform 1 0 384 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_98
timestamp 1626908933
transform 1 0 384 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_568
timestamp 1626908933
transform 1 0 960 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1198
timestamp 1626908933
transform 1 0 960 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_196
timestamp 1626908933
transform 1 0 1008 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_984
timestamp 1626908933
transform 1 0 1008 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_194
timestamp 1626908933
transform 1 0 1104 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_982
timestamp 1626908933
transform 1 0 1104 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_152
timestamp 1626908933
transform 1 0 1008 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_920
timestamp 1626908933
transform 1 0 1008 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_295
timestamp 1626908933
transform 1 0 1200 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1063
timestamp 1626908933
transform 1 0 1200 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_361
timestamp 1626908933
transform 1 0 1200 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1149
timestamp 1626908933
transform 1 0 1200 0 1 15651
box -29 -23 29 23
use M2M3_PR  M2M3_PR_30
timestamp 1626908933
transform 1 0 1296 0 1 16141
box -33 -37 33 37
use M2M3_PR  M2M3_PR_89
timestamp 1626908933
transform 1 0 1296 0 1 16141
box -33 -37 33 37
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_30
timestamp 1626908933
transform 1 0 1056 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_10
timestamp 1626908933
transform 1 0 1056 0 1 15984
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1410
timestamp 1626908933
transform 1 0 1488 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_642
timestamp 1626908933
transform 1 0 1488 0 1 15873
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_726
timestamp 1626908933
transform 1 0 1536 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_96
timestamp 1626908933
transform 1 0 1536 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1147
timestamp 1626908933
transform 1 0 1680 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_359
timestamp 1626908933
transform 1 0 1680 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_977
timestamp 1626908933
transform 1 0 1872 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_189
timestamp 1626908933
transform 1 0 1872 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1122
timestamp 1626908933
transform 1 0 1632 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_553
timestamp 1626908933
transform 1 0 1632 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_95
timestamp 1626908933
transform 1 0 2016 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_725
timestamp 1626908933
transform 1 0 2016 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_287
timestamp 1626908933
transform 1 0 2064 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1055
timestamp 1626908933
transform 1 0 2064 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_352
timestamp 1626908933
transform 1 0 2160 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1140
timestamp 1626908933
transform 1 0 2160 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_555
timestamp 1626908933
transform 1 0 2112 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1125
timestamp 1626908933
transform 1 0 2112 0 1 15984
box -38 -49 806 715
use L1M1_PR  L1M1_PR_186
timestamp 1626908933
transform 1 0 2352 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_974
timestamp 1626908933
transform 1 0 2352 0 1 15651
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_258
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_528
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_258
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_528
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_258
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_528
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_275
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_563
timestamp 1626908933
transform 1 0 2600 0 1 15984
box -200 -142 200 178
use L1M1_PR  L1M1_PR_110
timestamp 1626908933
transform 1 0 3216 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_898
timestamp 1626908933
transform 1 0 3216 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_31
timestamp 1626908933
transform 1 0 2880 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_11
timestamp 1626908933
transform 1 0 2880 0 1 15984
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1179
timestamp 1626908933
transform 1 0 3504 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_391
timestamp 1626908933
transform 1 0 3504 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1086
timestamp 1626908933
transform 1 0 3504 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_318
timestamp 1626908933
transform 1 0 3504 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_863
timestamp 1626908933
transform 1 0 3696 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_95
timestamp 1626908933
transform 1 0 3696 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_968
timestamp 1626908933
transform 1 0 4080 0 1 15799
box -29 -23 29 23
use L1M1_PR  L1M1_PR_180
timestamp 1626908933
transform 1 0 4080 0 1 15799
box -29 -23 29 23
use M1M2_PR  M1M2_PR_911
timestamp 1626908933
transform 1 0 4080 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_143
timestamp 1626908933
transform 1 0 4080 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_142
timestamp 1626908933
transform 1 0 4080 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_910
timestamp 1626908933
transform 1 0 4080 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_179
timestamp 1626908933
transform 1 0 4080 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_741
timestamp 1626908933
transform 1 0 3792 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_967
timestamp 1626908933
transform 1 0 4080 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1529
timestamp 1626908933
transform 1 0 3792 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_94
timestamp 1626908933
transform 1 0 3696 0 1 16243
box -32 -32 32 32
use M1M2_PR  M1M2_PR_862
timestamp 1626908933
transform 1 0 3696 0 1 16243
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_54
timestamp 1626908933
transform 1 0 3360 0 1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_134
timestamp 1626908933
transform 1 0 3360 0 1 15984
box -38 -49 902 715
use M1M2_PR  M1M2_PR_92
timestamp 1626908933
transform 1 0 4272 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_860
timestamp 1626908933
transform 1 0 4272 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_107
timestamp 1626908933
transform 1 0 4368 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_895
timestamp 1626908933
transform 1 0 4368 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_62
timestamp 1626908933
transform 1 0 4992 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_321
timestamp 1626908933
transform 1 0 4992 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_66
timestamp 1626908933
transform 1 0 5088 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_434
timestamp 1626908933
transform 1 0 5088 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_531
timestamp 1626908933
transform 1 0 4224 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1101
timestamp 1626908933
transform 1 0 4224 0 1 15984
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1519
timestamp 1626908933
transform 1 0 5136 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_751
timestamp 1626908933
transform 1 0 5136 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1563
timestamp 1626908933
transform 1 0 5232 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_886
timestamp 1626908933
transform 1 0 5328 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_775
timestamp 1626908933
transform 1 0 5232 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_98
timestamp 1626908933
transform 1 0 5328 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_724
timestamp 1626908933
transform 1 0 5280 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_94
timestamp 1626908933
transform 1 0 5280 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1081
timestamp 1626908933
transform 1 0 5376 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_512
timestamp 1626908933
transform 1 0 5376 0 1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_740
timestamp 1626908933
transform 1 0 6000 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1508
timestamp 1626908933
transform 1 0 6000 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_774
timestamp 1626908933
transform 1 0 5808 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1562
timestamp 1626908933
transform 1 0 5808 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_38
timestamp 1626908933
transform 1 0 5760 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_18
timestamp 1626908933
transform 1 0 5760 0 1 15984
box -38 -49 518 715
use L1M1_PR  L1M1_PR_172
timestamp 1626908933
transform 1 0 6192 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_960
timestamp 1626908933
transform 1 0 6192 0 1 15651
box -29 -23 29 23
use M2M3_PR  M2M3_PR_14
timestamp 1626908933
transform 1 0 6096 0 1 15775
box -33 -37 33 37
use M2M3_PR  M2M3_PR_73
timestamp 1626908933
transform 1 0 6096 0 1 15775
box -33 -37 33 37
use osc_core_VIA5  osc_core_VIA5_243
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_513
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_243
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_513
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_243
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_513
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_259
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_547
timestamp 1626908933
transform 1 0 6600 0 1 15984
box -200 -142 200 178
use L1M1_PR  L1M1_PR_929
timestamp 1626908933
transform 1 0 6096 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_141
timestamp 1626908933
transform 1 0 6096 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_887
timestamp 1626908933
transform 1 0 6096 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_119
timestamp 1626908933
transform 1 0 6096 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1199
timestamp 1626908933
transform 1 0 6432 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_569
timestamp 1626908933
transform 1 0 6432 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_709
timestamp 1626908933
transform 1 0 6240 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_341
timestamp 1626908933
transform 1 0 6240 0 1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1548
timestamp 1626908933
transform 1 0 6768 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_760
timestamp 1626908933
transform 1 0 6768 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1500
timestamp 1626908933
transform 1 0 6768 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_732
timestamp 1626908933
transform 1 0 6768 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1499
timestamp 1626908933
transform 1 0 6864 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_731
timestamp 1626908933
transform 1 0 6864 0 1 16169
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1547
timestamp 1626908933
transform 1 0 6864 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_759
timestamp 1626908933
transform 1 0 6864 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1498
timestamp 1626908933
transform 1 0 6864 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_730
timestamp 1626908933
transform 1 0 6864 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_56
timestamp 1626908933
transform 1 0 6528 0 1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_136
timestamp 1626908933
transform 1 0 6528 0 1 15984
box -38 -49 902 715
use L1M1_PR  L1M1_PR_959
timestamp 1626908933
transform 1 0 7056 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_171
timestamp 1626908933
transform 1 0 7056 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_903
timestamp 1626908933
transform 1 0 7056 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_135
timestamp 1626908933
transform 1 0 7056 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_958
timestamp 1626908933
transform 1 0 7056 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_170
timestamp 1626908933
transform 1 0 7056 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_902
timestamp 1626908933
transform 1 0 7056 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_134
timestamp 1626908933
transform 1 0 7056 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_710
timestamp 1626908933
transform 1 0 7392 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_342
timestamp 1626908933
transform 1 0 7392 0 1 15984
box -38 -49 230 715
use L1M1_PR  L1M1_PR_169
timestamp 1626908933
transform 1 0 7536 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_957
timestamp 1626908933
transform 1 0 7536 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_39
timestamp 1626908933
transform 1 0 7584 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_19
timestamp 1626908933
transform 1 0 7584 0 1 15984
box -38 -49 518 715
use M3M4_PR  M3M4_PR_34
timestamp 1626908933
transform 1 0 8064 0 1 15775
box -38 -33 38 33
use M3M4_PR  M3M4_PR_13
timestamp 1626908933
transform 1 0 8064 0 1 15775
box -38 -33 38 33
use M2M3_PR  M2M3_PR_66
timestamp 1626908933
transform 1 0 8112 0 1 15775
box -33 -37 33 37
use M2M3_PR  M2M3_PR_7
timestamp 1626908933
transform 1 0 8112 0 1 15775
box -33 -37 33 37
use M1M2_PR  M1M2_PR_877
timestamp 1626908933
transform 1 0 8112 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_109
timestamp 1626908933
transform 1 0 8112 0 1 15799
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1200
timestamp 1626908933
transform 1 0 8064 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_570
timestamp 1626908933
transform 1 0 8064 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1173
timestamp 1626908933
transform 1 0 8304 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_385
timestamp 1626908933
transform 1 0 8304 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1081
timestamp 1626908933
transform 1 0 8304 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_313
timestamp 1626908933
transform 1 0 8304 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_724
timestamp 1626908933
transform 1 0 8592 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1492
timestamp 1626908933
transform 1 0 8592 0 1 15799
box -32 -32 32 32
use L1M1_PR  L1M1_PR_128
timestamp 1626908933
transform 1 0 8496 0 1 15799
box -29 -23 29 23
use L1M1_PR  L1M1_PR_916
timestamp 1626908933
transform 1 0 8496 0 1 15799
box -29 -23 29 23
use M1M2_PR  M1M2_PR_723
timestamp 1626908933
transform 1 0 8592 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1491
timestamp 1626908933
transform 1 0 8592 0 1 16169
box -32 -32 32 32
use L1M1_PR  L1M1_PR_755
timestamp 1626908933
transform 1 0 8400 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1543
timestamp 1626908933
transform 1 0 8400 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_43
timestamp 1626908933
transform 1 0 8160 0 1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_123
timestamp 1626908933
transform 1 0 8160 0 1 15984
box -38 -49 902 715
use L1M1_PR  L1M1_PR_879
timestamp 1626908933
transform 1 0 8880 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_91
timestamp 1626908933
transform 1 0 8880 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_848
timestamp 1626908933
transform 1 0 8880 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_80
timestamp 1626908933
transform 1 0 8880 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_956
timestamp 1626908933
transform 1 0 8880 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_168
timestamp 1626908933
transform 1 0 8880 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_897
timestamp 1626908933
transform 1 0 8976 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_129
timestamp 1626908933
transform 1 0 8976 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1201
timestamp 1626908933
transform 1 0 9024 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_571
timestamp 1626908933
transform 1 0 9024 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1487
timestamp 1626908933
transform 1 0 9264 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_719
timestamp 1626908933
transform 1 0 9264 0 1 15873
box -32 -32 32 32
use L1M1_PR  L1M1_PR_744
timestamp 1626908933
transform 1 0 9552 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1532
timestamp 1626908933
transform 1 0 9552 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_90
timestamp 1626908933
transform 1 0 9648 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_733
timestamp 1626908933
transform 1 0 9360 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_878
timestamp 1626908933
transform 1 0 9648 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1521
timestamp 1626908933
transform 1 0 9360 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_37
timestamp 1626908933
transform 1 0 9120 0 1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_117
timestamp 1626908933
transform 1 0 9120 0 1 15984
box -38 -49 902 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_61
timestamp 1626908933
transform 1 0 9984 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_320
timestamp 1626908933
transform 1 0 9984 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_162
timestamp 1626908933
transform 1 0 9840 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_950
timestamp 1626908933
transform 1 0 9840 0 1 15651
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_228
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_498
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_228
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_498
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_228
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_498
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_243
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_531
timestamp 1626908933
transform 1 0 10600 0 1 15984
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_460
timestamp 1626908933
transform 1 0 10464 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1030
timestamp 1626908933
transform 1 0 10464 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_445
timestamp 1626908933
transform 1 0 10080 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1014
timestamp 1626908933
transform 1 0 10080 0 1 15984
box -38 -49 422 715
use L1M1_PR  L1M1_PR_158
timestamp 1626908933
transform 1 0 10896 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_742
timestamp 1626908933
transform 1 0 10608 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_946
timestamp 1626908933
transform 1 0 10896 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1530
timestamp 1626908933
transform 1 0 10608 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_700
timestamp 1626908933
transform 1 0 10896 0 1 15799
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1468
timestamp 1626908933
transform 1 0 10896 0 1 15799
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_572
timestamp 1626908933
transform 1 0 11232 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1202
timestamp 1626908933
transform 1 0 11232 0 1 15984
box -38 -49 134 715
use M2M3_PR  M2M3_PR_29
timestamp 1626908933
transform 1 0 11184 0 1 15775
box -33 -37 33 37
use M2M3_PR  M2M3_PR_88
timestamp 1626908933
transform 1 0 11184 0 1 15775
box -33 -37 33 37
use L1M1_PR  L1M1_PR_85
timestamp 1626908933
transform 1 0 11376 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_873
timestamp 1626908933
transform 1 0 11376 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_32
timestamp 1626908933
transform 1 0 11328 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_12
timestamp 1626908933
transform 1 0 11328 0 1 15984
box -38 -49 518 715
use M1M2_PR  M1M2_PR_128
timestamp 1626908933
transform 1 0 11664 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_896
timestamp 1626908933
transform 1 0 11664 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_65
timestamp 1626908933
transform 1 0 11808 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_433
timestamp 1626908933
transform 1 0 11808 0 1 15984
box -38 -49 230 715
use M1M2_PR  M1M2_PR_69
timestamp 1626908933
transform 1 0 12240 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_690
timestamp 1626908933
transform 1 0 11856 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_837
timestamp 1626908933
transform 1 0 12240 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1458
timestamp 1626908933
transform 1 0 11856 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_723
timestamp 1626908933
transform 1 0 11856 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1511
timestamp 1626908933
transform 1 0 11856 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_68
timestamp 1626908933
transform 1 0 12240 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_836
timestamp 1626908933
transform 1 0 12240 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_416
timestamp 1626908933
transform 1 0 12000 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_985
timestamp 1626908933
transform 1 0 12000 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1009
timestamp 1626908933
transform 1 0 12384 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_439
timestamp 1626908933
transform 1 0 12384 0 1 15984
box -38 -49 806 715
use L1M1_PR  L1M1_PR_869
timestamp 1626908933
transform 1 0 12240 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_81
timestamp 1626908933
transform 1 0 12240 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_13
timestamp 1626908933
transform 1 0 13152 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_33
timestamp 1626908933
transform 1 0 13152 0 1 15984
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1172
timestamp 1626908933
transform 1 0 13488 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_384
timestamp 1626908933
transform 1 0 13488 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1080
timestamp 1626908933
transform 1 0 13488 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_312
timestamp 1626908933
transform 1 0 13488 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_787
timestamp 1626908933
transform 1 0 13680 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_19
timestamp 1626908933
transform 1 0 13680 0 1 15651
box -32 -32 32 32
use osc_core_VIA3  osc_core_VIA3_5
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -28 96 28
use osc_core_VIA3  osc_core_VIA3_0
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_5
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -28 96 28
use osc_core_VIA2  osc_core_VIA2_0
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -28 96 28
use osc_core_VIA1  osc_core_VIA1_5
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -33 96 33
use osc_core_VIA1  osc_core_VIA1_0
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_5
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -33 96 33
use osc_core_VIA0  osc_core_VIA0_0
timestamp 1626908933
transform 1 0 14116 0 1 15802
box -97 -33 96 33
use M1M2_PR  M1M2_PR_18
timestamp 1626908933
transform 1 0 13680 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_786
timestamp 1626908933
transform 1 0 13680 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_14
timestamp 1626908933
transform 1 0 13488 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_802
timestamp 1626908933
transform 1 0 13488 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_423
timestamp 1626908933
transform 1 0 13632 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_993
timestamp 1626908933
transform 1 0 13632 0 1 15984
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_515
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_227
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -142 200 178
use L1M1_PR  L1M1_PR_800
timestamp 1626908933
transform 1 0 14448 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_12
timestamp 1626908933
transform 1 0 14448 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_784
timestamp 1626908933
transform 1 0 14544 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_16
timestamp 1626908933
transform 1 0 14544 0 1 15651
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_483
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_213
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_483
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_213
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_483
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_213
timestamp 1626908933
transform 1 0 14600 0 1 15984
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_60
timestamp 1626908933
transform 1 0 14976 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_319
timestamp 1626908933
transform 1 0 14976 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_343
timestamp 1626908933
transform 1 0 14784 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_711
timestamp 1626908933
transform 1 0 14784 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_369
timestamp 1626908933
transform 1 0 14400 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_938
timestamp 1626908933
transform 1 0 14400 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_432
timestamp 1626908933
transform 1 0 15072 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_64
timestamp 1626908933
transform 1 0 15072 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_954
timestamp 1626908933
transform 1 0 15264 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_384
timestamp 1626908933
transform 1 0 15264 0 1 15984
box -38 -49 806 715
use M2M3_PR  M2M3_PR_62
timestamp 1626908933
transform 1 0 15312 0 1 15897
box -33 -37 33 37
use M2M3_PR  M2M3_PR_3
timestamp 1626908933
transform 1 0 15312 0 1 15897
box -33 -37 33 37
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_16
timestamp 1626908933
transform 1 0 16032 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_36
timestamp 1626908933
transform 1 0 16032 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_928
timestamp 1626908933
transform 1 0 16704 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_358
timestamp 1626908933
transform 1 0 16704 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_431
timestamp 1626908933
transform 1 0 16512 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_63
timestamp 1626908933
transform 1 0 16512 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_712
timestamp 1626908933
transform 1 0 17568 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_344
timestamp 1626908933
transform 1 0 17568 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_318
timestamp 1626908933
transform 1 0 17472 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_59
timestamp 1626908933
transform 1 0 17472 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1203
timestamp 1626908933
transform 1 0 17760 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_573
timestamp 1626908933
transform 1 0 17760 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_908
timestamp 1626908933
transform 1 0 17808 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_120
timestamp 1626908933
transform 1 0 17808 0 1 16095
box -29 -23 29 23
use M1M2_PR  M1M2_PR_872
timestamp 1626908933
transform 1 0 17808 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_104
timestamp 1626908933
transform 1 0 17808 0 1 16095
box -32 -32 32 32
use M3M4_PR  M3M4_PR_24
timestamp 1626908933
transform 1 0 17904 0 1 15897
box -38 -33 38 33
use M3M4_PR  M3M4_PR_3
timestamp 1626908933
transform 1 0 17904 0 1 15897
box -38 -33 38 33
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_17
timestamp 1626908933
transform 1 0 17856 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_37
timestamp 1626908933
transform 1 0 17856 0 1 15984
box -38 -49 518 715
use M1M2_PR  M1M2_PR_776
timestamp 1626908933
transform 1 0 18096 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_8
timestamp 1626908933
transform 1 0 18096 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_777
timestamp 1626908933
transform 1 0 18096 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_9
timestamp 1626908933
transform 1 0 18096 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1408
timestamp 1626908933
transform 1 0 18288 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_620
timestamp 1626908933
transform 1 0 18288 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1312
timestamp 1626908933
transform 1 0 18288 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_544
timestamp 1626908933
transform 1 0 18288 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_723
timestamp 1626908933
transform 1 0 18336 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_93
timestamp 1626908933
transform 1 0 18336 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_907
timestamp 1626908933
transform 1 0 18768 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_119
timestamp 1626908933
transform 1 0 18768 0 1 15651
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_499
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_211
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_468
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_198
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_468
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_198
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_468
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_198
timestamp 1626908933
transform 1 0 18600 0 1 15984
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_295
timestamp 1626908933
transform 1 0 18432 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_864
timestamp 1626908933
transform 1 0 18432 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_335
timestamp 1626908933
transform 1 0 18816 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_905
timestamp 1626908933
transform 1 0 18816 0 1 15984
box -38 -49 806 715
use M1M2_PR  M1M2_PR_775
timestamp 1626908933
transform 1 0 19536 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_7
timestamp 1626908933
transform 1 0 19536 0 1 16169
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_848
timestamp 1626908933
transform 1 0 19584 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_279
timestamp 1626908933
transform 1 0 19584 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_14
timestamp 1626908933
transform 1 0 20160 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_34
timestamp 1626908933
transform 1 0 20160 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1204
timestamp 1626908933
transform 1 0 20064 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_574
timestamp 1626908933
transform 1 0 20064 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_317
timestamp 1626908933
transform 1 0 19968 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_58
timestamp 1626908933
transform 1 0 19968 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_855
timestamp 1626908933
transform 1 0 20736 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_285
timestamp 1626908933
transform 1 0 20736 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_722
timestamp 1626908933
transform 1 0 20640 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_92
timestamp 1626908933
transform 1 0 20640 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_815
timestamp 1626908933
transform 1 0 21504 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_246
timestamp 1626908933
transform 1 0 21504 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_91
timestamp 1626908933
transform 1 0 21888 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_721
timestamp 1626908933
transform 1 0 21888 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_550
timestamp 1626908933
transform 1 0 21936 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1318
timestamp 1626908933
transform 1 0 21936 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_626
timestamp 1626908933
transform 1 0 21936 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1414
timestamp 1626908933
transform 1 0 21936 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_549
timestamp 1626908933
transform 1 0 21936 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1317
timestamp 1626908933
transform 1 0 21936 0 1 16095
box -32 -32 32 32
use M1M2_PR  M1M2_PR_810
timestamp 1626908933
transform 1 0 22320 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_42
timestamp 1626908933
transform 1 0 22320 0 1 15651
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_483
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_195
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -142 200 178
use M1M2_PR  M1M2_PR_773
timestamp 1626908933
transform 1 0 22128 0 1 16169
box -32 -32 32 32
use M1M2_PR  M1M2_PR_5
timestamp 1626908933
transform 1 0 22128 0 1 16169
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_453
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_183
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_453
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_183
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_453
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_183
timestamp 1626908933
transform 1 0 22600 0 1 15984
box -200 -49 200 49
use L1M1_PR  L1M1_PR_833
timestamp 1626908933
transform 1 0 22320 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_45
timestamp 1626908933
transform 1 0 22320 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_809
timestamp 1626908933
transform 1 0 22320 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_41
timestamp 1626908933
transform 1 0 22320 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_35
timestamp 1626908933
transform 1 0 21984 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_15
timestamp 1626908933
transform 1 0 21984 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_57
timestamp 1626908933
transform 1 0 22464 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_316
timestamp 1626908933
transform 1 0 22464 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_90
timestamp 1626908933
transform 1 0 22560 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_720
timestamp 1626908933
transform 1 0 22560 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_44
timestamp 1626908933
transform 1 0 22800 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_832
timestamp 1626908933
transform 1 0 22800 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_36
timestamp 1626908933
transform 1 0 22992 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_804
timestamp 1626908933
transform 1 0 22992 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_247
timestamp 1626908933
transform 1 0 22656 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_817
timestamp 1626908933
transform 1 0 22656 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_783
timestamp 1626908933
transform 1 0 23424 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_214
timestamp 1626908933
transform 1 0 23424 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_89
timestamp 1626908933
transform 1 0 23808 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_719
timestamp 1626908933
transform 1 0 23808 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1196
timestamp 1626908933
transform 1 0 24048 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_428
timestamp 1626908933
transform 1 0 24048 0 1 15651
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1282
timestamp 1626908933
transform 1 0 24336 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_494
timestamp 1626908933
transform 1 0 24336 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1219
timestamp 1626908933
transform 1 0 24336 0 1 15799
box -29 -23 29 23
use L1M1_PR  L1M1_PR_431
timestamp 1626908933
transform 1 0 24336 0 1 15799
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1413
timestamp 1626908933
transform 1 0 24048 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_625
timestamp 1626908933
transform 1 0 24048 0 1 16095
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1221
timestamp 1626908933
transform 1 0 24240 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_433
timestamp 1626908933
transform 1 0 24240 0 1 16317
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1128
timestamp 1626908933
transform 1 0 24144 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_360
timestamp 1626908933
transform 1 0 24144 0 1 16317
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1218
timestamp 1626908933
transform 1 0 24336 0 1 16317
box -29 -23 29 23
use L1M1_PR  L1M1_PR_430
timestamp 1626908933
transform 1 0 24336 0 1 16317
box -29 -23 29 23
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_1
timestamp 1626908933
transform -1 0 24384 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_3
timestamp 1626908933
transform -1 0 24384 0 1 15984
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_88
timestamp 1626908933
transform 1 0 24384 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_718
timestamp 1626908933
transform 1 0 24384 0 1 15984
box -38 -49 134 715
use M1M2_PR  M1M2_PR_359
timestamp 1626908933
transform 1 0 24528 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1127
timestamp 1626908933
transform 1 0 24528 0 1 15873
box -32 -32 32 32
use M1M2_PR  M1M2_PR_358
timestamp 1626908933
transform 1 0 24528 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1126
timestamp 1626908933
transform 1 0 24528 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_315
timestamp 1626908933
transform 1 0 24960 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_56
timestamp 1626908933
transform 1 0 24960 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1290
timestamp 1626908933
transform 1 0 24912 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_502
timestamp 1626908933
transform 1 0 24912 0 1 15651
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_717
timestamp 1626908933
transform 1 0 24864 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_87
timestamp 1626908933
transform 1 0 24864 0 1 15984
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1297
timestamp 1626908933
transform 1 0 25200 0 1 15651
box -29 -23 29 23
use L1M1_PR  L1M1_PR_509
timestamp 1626908933
transform 1 0 25200 0 1 15651
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1220
timestamp 1626908933
transform 1 0 25200 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_452
timestamp 1626908933
transform 1 0 25200 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_430
timestamp 1626908933
transform 1 0 25056 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_62
timestamp 1626908933
transform 1 0 25056 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_208
timestamp 1626908933
transform 1 0 24480 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_777
timestamp 1626908933
transform 1 0 24480 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_775
timestamp 1626908933
transform 1 0 25248 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_205
timestamp 1626908933
transform 1 0 25248 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_747
timestamp 1626908933
transform 1 0 26016 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_178
timestamp 1626908933
transform 1 0 26016 0 1 15984
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_467
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_179
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_438
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_168
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_438
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_168
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_438
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_168
timestamp 1626908933
transform 1 0 26600 0 1 15984
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_716
timestamp 1626908933
transform 1 0 26400 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_86
timestamp 1626908933
transform 1 0 26400 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_183
timestamp 1626908933
transform 1 0 26496 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_753
timestamp 1626908933
transform 1 0 26496 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_61
timestamp 1626908933
transform 1 0 27552 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_429
timestamp 1626908933
transform 1 0 27552 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_55
timestamp 1626908933
transform 1 0 27456 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_314
timestamp 1626908933
transform 1 0 27456 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_575
timestamp 1626908933
transform 1 0 27360 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1205
timestamp 1626908933
transform 1 0 27360 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_85
timestamp 1626908933
transform 1 0 27264 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_715
timestamp 1626908933
transform 1 0 27264 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_84
timestamp 1626908933
transform 1 0 27744 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_714
timestamp 1626908933
transform 1 0 27744 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_159
timestamp 1626908933
transform 1 0 27840 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_729
timestamp 1626908933
transform 1 0 27840 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_710
timestamp 1626908933
transform 1 0 28608 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_141
timestamp 1626908933
transform 1 0 28608 0 1 15984
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1191
timestamp 1626908933
transform 1 0 29040 0 1 15651
box -32 -32 32 32
use M1M2_PR  M1M2_PR_423
timestamp 1626908933
transform 1 0 29040 0 1 15651
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_713
timestamp 1626908933
transform 1 0 28992 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_83
timestamp 1626908933
transform 1 0 28992 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_705
timestamp 1626908933
transform 1 0 29088 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_135
timestamp 1626908933
transform 1 0 29088 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1206
timestamp 1626908933
transform 1 0 29856 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_576
timestamp 1626908933
transform 1 0 29856 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_82
timestamp 1626908933
transform 1 0 30240 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_712
timestamp 1626908933
transform 1 0 30240 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_60
timestamp 1626908933
transform 1 0 30048 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_428
timestamp 1626908933
transform 1 0 30048 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_54
timestamp 1626908933
transform 1 0 29952 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_313
timestamp 1626908933
transform 1 0 29952 0 1 15984
box -38 -49 134 715
use osc_core_VIA5  osc_core_VIA5_153
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_423
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_153
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_423
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_153
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_423
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_163
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_451
timestamp 1626908933
transform 1 0 30600 0 1 15984
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_110
timestamp 1626908933
transform 1 0 30336 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_680
timestamp 1626908933
transform 1 0 30336 0 1 15984
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1374
timestamp 1626908933
transform 1 0 30960 0 1 16317
box -32 -32 32 32
use M1M2_PR  M1M2_PR_606
timestamp 1626908933
transform 1 0 30960 0 1 16317
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_427
timestamp 1626908933
transform 1 0 31104 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_59
timestamp 1626908933
transform 1 0 31104 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_658
timestamp 1626908933
transform 1 0 31296 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_89
timestamp 1626908933
transform 1 0 31296 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_650
timestamp 1626908933
transform 1 0 31680 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_80
timestamp 1626908933
transform 1 0 31680 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_625
timestamp 1626908933
transform 1 0 32544 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_56
timestamp 1626908933
transform 1 0 32544 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_711
timestamp 1626908933
transform 1 0 32448 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_81
timestamp 1626908933
transform 1 0 32448 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_620
timestamp 1626908933
transform 1 0 32928 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_50
timestamp 1626908933
transform 1 0 32928 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_710
timestamp 1626908933
transform 1 0 33696 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_80
timestamp 1626908933
transform 1 0 33696 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_592
timestamp 1626908933
transform 1 0 33792 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_23
timestamp 1626908933
transform 1 0 33792 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_590
timestamp 1626908933
transform 1 0 34176 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_20
timestamp 1626908933
transform 1 0 34176 0 1 15984
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_408
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_138
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_408
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_138
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_408
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_138
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_147
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_435
timestamp 1626908933
transform 1 0 34600 0 1 15984
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_53
timestamp 1626908933
transform 1 0 34944 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_312
timestamp 1626908933
transform 1 0 34944 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_345
timestamp 1626908933
transform 1 0 35424 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_713
timestamp 1626908933
transform 1 0 35424 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_577
timestamp 1626908933
transform 1 0 35616 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1207
timestamp 1626908933
transform 1 0 35616 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_3
timestamp 1626908933
transform 1 0 35040 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_572
timestamp 1626908933
transform 1 0 35040 0 1 15984
box -38 -49 422 715
use M2M3_PR_R  M2M3_PR_R_3
timestamp 1626908933
transform 1 0 48 0 1 17117
box -37 -33 37 33
use M2M3_PR_R  M2M3_PR_R_1
timestamp 1626908933
transform 1 0 48 0 1 17117
box -37 -33 37 33
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1138
timestamp 1626908933
transform 1 0 288 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_568
timestamp 1626908933
transform 1 0 288 0 -1 17316
box -38 -49 806 715
use M2M3_PR  M2M3_PR_104
timestamp 1626908933
transform 1 0 48 0 1 16507
box -33 -37 33 37
use M2M3_PR  M2M3_PR_45
timestamp 1626908933
transform 1 0 48 0 1 16507
box -33 -37 33 37
use osc_core_VIA4  osc_core_VIA4_131
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_419
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_392
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_122
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_392
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_122
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_392
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_122
timestamp 1626908933
transform 1 0 600 0 1 16650
box -200 -49 200 49
use M1M2_PR  M1M2_PR_934
timestamp 1626908933
transform 1 0 1104 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_166
timestamp 1626908933
transform 1 0 1104 0 1 16539
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_0
timestamp 1626908933
transform 1 0 1056 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_10
timestamp 1626908933
transform 1 0 1056 0 -1 17316
box -38 -49 518 715
use M1M2_PR  M1M2_PR_930
timestamp 1626908933
transform 1 0 1200 0 1 16835
box -32 -32 32 32
use M1M2_PR  M1M2_PR_162
timestamp 1626908933
transform 1 0 1200 0 1 16835
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1420
timestamp 1626908933
transform 1 0 1296 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_632
timestamp 1626908933
transform 1 0 1296 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1326
timestamp 1626908933
transform 1 0 1296 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_558
timestamp 1626908933
transform 1 0 1296 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_998
timestamp 1626908933
transform 1 0 1200 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_210
timestamp 1626908933
transform 1 0 1200 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_996
timestamp 1626908933
transform 1 0 1584 0 1 16835
box -29 -23 29 23
use L1M1_PR  L1M1_PR_208
timestamp 1626908933
transform 1 0 1584 0 1 16835
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1124
timestamp 1626908933
transform 1 0 1728 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_554
timestamp 1626908933
transform 1 0 1728 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_426
timestamp 1626908933
transform 1 0 1536 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_58
timestamp 1626908933
transform 1 0 1536 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_346
timestamp 1626908933
transform 1 0 2592 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_714
timestamp 1626908933
transform 1 0 2592 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_578
timestamp 1626908933
transform 1 0 2784 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1208
timestamp 1626908933
transform 1 0 2784 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_52
timestamp 1626908933
transform 1 0 2496 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_311
timestamp 1626908933
transform 1 0 2496 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_939
timestamp 1626908933
transform 1 0 2928 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_171
timestamp 1626908933
transform 1 0 2928 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1003
timestamp 1626908933
transform 1 0 3024 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_215
timestamp 1626908933
transform 1 0 3024 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_935
timestamp 1626908933
transform 1 0 3024 0 1 16835
box -32 -32 32 32
use M1M2_PR  M1M2_PR_167
timestamp 1626908933
transform 1 0 3024 0 1 16835
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1424
timestamp 1626908933
transform 1 0 3120 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_636
timestamp 1626908933
transform 1 0 3120 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1339
timestamp 1626908933
transform 1 0 3120 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_571
timestamp 1626908933
transform 1 0 3120 0 1 16983
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_1
timestamp 1626908933
transform 1 0 2880 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_11
timestamp 1626908933
transform 1 0 2880 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_347
timestamp 1626908933
transform 1 0 3360 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_715
timestamp 1626908933
transform 1 0 3360 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_579
timestamp 1626908933
transform 1 0 3552 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1209
timestamp 1626908933
transform 1 0 3552 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_213
timestamp 1626908933
transform 1 0 3408 0 1 16835
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1001
timestamp 1626908933
transform 1 0 3408 0 1 16835
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1482
timestamp 1626908933
transform 1 0 3792 0 1 16465
box -32 -32 32 32
use M1M2_PR  M1M2_PR_714
timestamp 1626908933
transform 1 0 3792 0 1 16465
box -32 -32 32 32
use M2M3_PR  M2M3_PR_115
timestamp 1626908933
transform 1 0 3792 0 1 16873
box -33 -37 33 37
use M2M3_PR  M2M3_PR_56
timestamp 1626908933
transform 1 0 3792 0 1 16873
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1481
timestamp 1626908933
transform 1 0 3792 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_713
timestamp 1626908933
transform 1 0 3792 0 1 16909
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1528
timestamp 1626908933
transform 1 0 3888 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_740
timestamp 1626908933
transform 1 0 3888 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_861
timestamp 1626908933
transform 1 0 3984 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_93
timestamp 1626908933
transform 1 0 3984 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_909
timestamp 1626908933
transform 1 0 4176 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_141
timestamp 1626908933
transform 1 0 4176 0 1 16983
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_55
timestamp 1626908933
transform 1 0 3648 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_135
timestamp 1626908933
transform 1 0 3648 0 -1 17316
box -38 -49 902 715
use osc_core_VIA5  osc_core_VIA5_107
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_377
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_107
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_377
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_107
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_377
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_115
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_403
timestamp 1626908933
transform 1 0 4600 0 1 16650
box -200 -142 200 178
use L1M1_PR  L1M1_PR_966
timestamp 1626908933
transform 1 0 4176 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_178
timestamp 1626908933
transform 1 0 4176 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_891
timestamp 1626908933
transform 1 0 4656 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_103
timestamp 1626908933
transform 1 0 4656 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1565
timestamp 1626908933
transform 1 0 4944 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_777
timestamp 1626908933
transform 1 0 4944 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1520
timestamp 1626908933
transform 1 0 4944 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1396
timestamp 1626908933
transform 1 0 5040 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_752
timestamp 1626908933
transform 1 0 4944 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_628
timestamp 1626908933
transform 1 0 5040 0 1 16983
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_46
timestamp 1626908933
transform -1 0 5376 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_126
timestamp 1626908933
transform -1 0 5376 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_511
timestamp 1626908933
transform 1 0 5376 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1080
timestamp 1626908933
transform 1 0 5376 0 -1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_230
timestamp 1626908933
transform 1 0 5904 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_234
timestamp 1626908933
transform 1 0 5808 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_998
timestamp 1626908933
transform 1 0 5904 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1002
timestamp 1626908933
transform 1 0 5808 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_285
timestamp 1626908933
transform 1 0 5904 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1073
timestamp 1626908933
transform 1 0 5904 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_664
timestamp 1626908933
transform 1 0 5904 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1452
timestamp 1626908933
transform 1 0 5904 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_8
timestamp 1626908933
transform 1 0 5760 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_18
timestamp 1626908933
transform 1 0 5760 0 -1 17316
box -38 -49 518 715
use M1M2_PR  M1M2_PR_1404
timestamp 1626908933
transform 1 0 6864 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_636
timestamp 1626908933
transform 1 0 6864 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1072
timestamp 1626908933
transform 1 0 6288 0 1 16761
box -29 -23 29 23
use L1M1_PR  L1M1_PR_284
timestamp 1626908933
transform 1 0 6288 0 1 16761
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_10
timestamp 1626908933
transform 1 0 6240 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_1
timestamp 1626908933
transform 1 0 6240 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1075
timestamp 1626908933
transform 1 0 6624 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_505
timestamp 1626908933
transform 1 0 6624 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_580
timestamp 1626908933
transform 1 0 7392 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1210
timestamp 1626908933
transform 1 0 7392 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_310
timestamp 1626908933
transform 1 0 7488 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_51
timestamp 1626908933
transform 1 0 7488 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1456
timestamp 1626908933
transform 1 0 7728 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_668
timestamp 1626908933
transform 1 0 7728 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1006
timestamp 1626908933
transform 1 0 7632 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_238
timestamp 1626908933
transform 1 0 7632 0 1 17057
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1079
timestamp 1626908933
transform 1 0 7728 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_291
timestamp 1626908933
transform 1 0 7728 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1007
timestamp 1626908933
transform 1 0 7632 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_239
timestamp 1626908933
transform 1 0 7632 0 1 16539
box -32 -32 32 32
use M2M3_PR  M2M3_PR_103
timestamp 1626908933
transform 1 0 7824 0 1 16507
box -33 -37 33 37
use M2M3_PR  M2M3_PR_44
timestamp 1626908933
transform 1 0 7824 0 1 16507
box -33 -37 33 37
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_9
timestamp 1626908933
transform 1 0 7584 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_19
timestamp 1626908933
transform 1 0 7584 0 -1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1077
timestamp 1626908933
transform 1 0 8016 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_289
timestamp 1626908933
transform 1 0 8016 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1211
timestamp 1626908933
transform 1 0 8064 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_581
timestamp 1626908933
transform 1 0 8064 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_704
timestamp 1626908933
transform 1 0 8304 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1472
timestamp 1626908933
transform 1 0 8304 0 1 16539
box -32 -32 32 32
use M2M3_PR  M2M3_PR_55
timestamp 1626908933
transform 1 0 8304 0 1 16873
box -33 -37 33 37
use M2M3_PR  M2M3_PR_114
timestamp 1626908933
transform 1 0 8304 0 1 16873
box -33 -37 33 37
use M1M2_PR  M1M2_PR_703
timestamp 1626908933
transform 1 0 8304 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1471
timestamp 1626908933
transform 1 0 8304 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_736
timestamp 1626908933
transform 1 0 8304 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1524
timestamp 1626908933
transform 1 0 8304 0 1 16983
box -29 -23 29 23
use M2M3_PR  M2M3_PR_43
timestamp 1626908933
transform 1 0 8304 0 1 17117
box -33 -37 33 37
use M2M3_PR  M2M3_PR_102
timestamp 1626908933
transform 1 0 8304 0 1 17117
box -33 -37 33 37
use osc_core_VIA7  osc_core_VIA7_362
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_92
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_362
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_92
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_362
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_92
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_387
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_99
timestamp 1626908933
transform 1 0 8600 0 1 16650
box -200 -142 200 178
use L1M1_PR  L1M1_PR_880
timestamp 1626908933
transform 1 0 8688 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_92
timestamp 1626908933
transform 1 0 8688 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_38
timestamp 1626908933
transform 1 0 8160 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_118
timestamp 1626908933
transform 1 0 8160 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_348
timestamp 1626908933
transform 1 0 9024 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_716
timestamp 1626908933
transform 1 0 9024 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_79
timestamp 1626908933
transform 1 0 8880 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_718
timestamp 1626908933
transform 1 0 9264 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_847
timestamp 1626908933
transform 1 0 8880 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1486
timestamp 1626908933
transform 1 0 9264 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_78
timestamp 1626908933
transform 1 0 9648 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_846
timestamp 1626908933
transform 1 0 9648 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_746
timestamp 1626908933
transform 1 0 9360 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1534
timestamp 1626908933
transform 1 0 9360 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_41
timestamp 1626908933
transform 1 0 9216 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_121
timestamp 1626908933
transform 1 0 9216 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_349
timestamp 1626908933
transform 1 0 10080 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_717
timestamp 1626908933
transform 1 0 10080 0 -1 17316
box -38 -49 230 715
use L1M1_PR  L1M1_PR_87
timestamp 1626908933
transform 1 0 9744 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_875
timestamp 1626908933
transform 1 0 9744 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_582
timestamp 1626908933
transform 1 0 10272 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1212
timestamp 1626908933
transform 1 0 10272 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_702
timestamp 1626908933
transform 1 0 10512 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1470
timestamp 1626908933
transform 1 0 10512 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_701
timestamp 1626908933
transform 1 0 10512 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1469
timestamp 1626908933
transform 1 0 10512 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_731
timestamp 1626908933
transform 1 0 10512 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1519
timestamp 1626908933
transform 1 0 10512 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_39
timestamp 1626908933
transform 1 0 10368 0 -1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_119
timestamp 1626908933
transform 1 0 10368 0 -1 17316
box -38 -49 902 715
use L1M1_PR  L1M1_PR_86
timestamp 1626908933
transform 1 0 10896 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_874
timestamp 1626908933
transform 1 0 10896 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1213
timestamp 1626908933
transform 1 0 11232 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_583
timestamp 1626908933
transform 1 0 11232 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_951
timestamp 1626908933
transform 1 0 11376 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_183
timestamp 1626908933
transform 1 0 11376 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_947
timestamp 1626908933
transform 1 0 11568 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_179
timestamp 1626908933
transform 1 0 11568 0 1 16983
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1428
timestamp 1626908933
transform 1 0 11472 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_640
timestamp 1626908933
transform 1 0 11472 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1016
timestamp 1626908933
transform 1 0 11472 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_228
timestamp 1626908933
transform 1 0 11472 0 1 16539
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_2
timestamp 1626908933
transform 1 0 11328 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_12
timestamp 1626908933
transform 1 0 11328 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_79
timestamp 1626908933
transform 1 0 12000 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_709
timestamp 1626908933
transform 1 0 12000 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_57
timestamp 1626908933
transform 1 0 11808 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_425
timestamp 1626908933
transform 1 0 11808 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_127
timestamp 1626908933
transform 1 0 11664 0 1 16465
box -32 -32 32 32
use M1M2_PR  M1M2_PR_895
timestamp 1626908933
transform 1 0 11664 0 1 16465
box -32 -32 32 32
use L1M1_PR  L1M1_PR_227
timestamp 1626908933
transform 1 0 11760 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1015
timestamp 1626908933
transform 1 0 11760 0 1 16983
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_371
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_83
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_347
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_77
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_347
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_77
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_347
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_77
timestamp 1626908933
transform 1 0 12600 0 1 16650
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_984
timestamp 1626908933
transform 1 0 12096 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_415
timestamp 1626908933
transform 1 0 12096 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_50
timestamp 1626908933
transform 1 0 12480 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_309
timestamp 1626908933
transform 1 0 12480 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_56
timestamp 1626908933
transform 1 0 12576 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_424
timestamp 1626908933
transform 1 0 12576 0 -1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_188
timestamp 1626908933
transform 1 0 13104 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_956
timestamp 1626908933
transform 1 0 13104 0 1 16539
box -32 -32 32 32
use L1M1_PR  L1M1_PR_234
timestamp 1626908933
transform 1 0 13296 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1022
timestamp 1626908933
transform 1 0 13296 0 1 16539
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_3
timestamp 1626908933
transform 1 0 13152 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_13
timestamp 1626908933
transform 1 0 13152 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_391
timestamp 1626908933
transform 1 0 12768 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_960
timestamp 1626908933
transform 1 0 12768 0 -1 17316
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1432
timestamp 1626908933
transform 1 0 13392 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_644
timestamp 1626908933
transform 1 0 13392 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_2
timestamp 1626908933
transform 1 0 13632 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_0
timestamp 1626908933
transform 1 0 13632 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_937
timestamp 1626908933
transform 1 0 14400 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_368
timestamp 1626908933
transform 1 0 14400 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_423
timestamp 1626908933
transform 1 0 14784 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_55
timestamp 1626908933
transform 1 0 14784 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_975
timestamp 1626908933
transform 1 0 14976 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_405
timestamp 1626908933
transform 1 0 14976 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_54
timestamp 1626908933
transform 1 0 15744 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_422
timestamp 1626908933
transform 1 0 15744 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_584
timestamp 1626908933
transform 1 0 15936 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1214
timestamp 1626908933
transform 1 0 15936 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_156
timestamp 1626908933
transform 1 0 15984 0 1 16465
box -29 -23 29 23
use L1M1_PR  L1M1_PR_944
timestamp 1626908933
transform 1 0 15984 0 1 16465
box -29 -23 29 23
use M1M2_PR  M1M2_PR_579
timestamp 1626908933
transform 1 0 15792 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1347
timestamp 1626908933
transform 1 0 15792 0 1 16983
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_6
timestamp 1626908933
transform 1 0 16032 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_16
timestamp 1626908933
transform 1 0 16032 0 -1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1055
timestamp 1626908933
transform 1 0 16176 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_267
timestamp 1626908933
transform 1 0 16176 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_986
timestamp 1626908933
transform 1 0 16272 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_218
timestamp 1626908933
transform 1 0 16272 0 1 16539
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_332
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_62
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_332
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_62
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_332
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_62
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_67
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_355
timestamp 1626908933
transform 1 0 16600 0 1 16650
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1444
timestamp 1626908933
transform 1 0 16272 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_656
timestamp 1626908933
transform 1 0 16272 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_981
timestamp 1626908933
transform 1 0 16464 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_213
timestamp 1626908933
transform 1 0 16464 0 1 17131
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_53
timestamp 1626908933
transform 1 0 16512 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_421
timestamp 1626908933
transform 1 0 16512 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_357
timestamp 1626908933
transform 1 0 16704 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_927
timestamp 1626908933
transform 1 0 16704 0 -1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_608
timestamp 1626908933
transform 1 0 17040 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1376
timestamp 1626908933
transform 1 0 17040 0 1 16391
box -32 -32 32 32
use M1M2_PR  M1M2_PR_607
timestamp 1626908933
transform 1 0 17040 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1375
timestamp 1626908933
transform 1 0 17040 0 1 17057
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_350
timestamp 1626908933
transform 1 0 17568 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_718
timestamp 1626908933
transform 1 0 17568 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_49
timestamp 1626908933
transform 1 0 17472 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_308
timestamp 1626908933
transform 1 0 17472 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_585
timestamp 1626908933
transform 1 0 17760 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1215
timestamp 1626908933
transform 1 0 17760 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_988
timestamp 1626908933
transform 1 0 17904 0 1 17057
box -32 -32 32 32
use M1M2_PR  M1M2_PR_220
timestamp 1626908933
transform 1 0 17904 0 1 17057
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_17
timestamp 1626908933
transform 1 0 17856 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_7
timestamp 1626908933
transform 1 0 17856 0 -1 17316
box -38 -49 518 715
use M1M2_PR  M1M2_PR_991
timestamp 1626908933
transform 1 0 17808 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_223
timestamp 1626908933
transform 1 0 17808 0 1 16539
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_78
timestamp 1626908933
transform 1 0 18336 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_708
timestamp 1626908933
transform 1 0 18336 0 -1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_272
timestamp 1626908933
transform 1 0 18000 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1060
timestamp 1626908933
transform 1 0 18000 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_270
timestamp 1626908933
transform 1 0 18288 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_660
timestamp 1626908933
transform 1 0 18000 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1058
timestamp 1626908933
transform 1 0 18288 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1448
timestamp 1626908933
transform 1 0 18000 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_334
timestamp 1626908933
transform 1 0 18816 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_904
timestamp 1626908933
transform 1 0 18816 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_294
timestamp 1626908933
transform 1 0 18432 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_863
timestamp 1626908933
transform 1 0 18432 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_847
timestamp 1626908933
transform 1 0 19584 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_278
timestamp 1626908933
transform 1 0 19584 0 -1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_774
timestamp 1626908933
transform 1 0 19536 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_6
timestamp 1626908933
transform 1 0 19536 0 1 16539
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_77
timestamp 1626908933
transform 1 0 19968 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_586
timestamp 1626908933
transform 1 0 20064 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_707
timestamp 1626908933
transform 1 0 19968 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1216
timestamp 1626908933
transform 1 0 20064 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_620
timestamp 1626908933
transform 1 0 19920 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1388
timestamp 1626908933
transform 1 0 19920 0 1 16909
box -32 -32 32 32
use L1M1_PR  L1M1_PR_793
timestamp 1626908933
transform 1 0 20112 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_5
timestamp 1626908933
transform 1 0 20112 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1036
timestamp 1626908933
transform 1 0 20304 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_248
timestamp 1626908933
transform 1 0 20304 0 1 16539
box -29 -23 29 23
use M1M2_PR  M1M2_PR_969
timestamp 1626908933
transform 1 0 20304 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_201
timestamp 1626908933
transform 1 0 20304 0 1 16539
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_317
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_47
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_317
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_47
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_317
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_47
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_339
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_51
timestamp 1626908933
transform 1 0 20600 0 1 16650
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1436
timestamp 1626908933
transform 1 0 20304 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_648
timestamp 1626908933
transform 1 0 20304 0 1 16983
box -29 -23 29 23
use M1M2_PR  M1M2_PR_966
timestamp 1626908933
transform 1 0 20400 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_198
timestamp 1626908933
transform 1 0 20400 0 1 16983
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_4
timestamp 1626908933
transform 1 0 20160 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_14
timestamp 1626908933
transform 1 0 20160 0 -1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1034
timestamp 1626908933
transform 1 0 20592 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_246
timestamp 1626908933
transform 1 0 20592 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_854
timestamp 1626908933
transform 1 0 20736 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_284
timestamp 1626908933
transform 1 0 20736 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_706
timestamp 1626908933
transform 1 0 20640 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_76
timestamp 1626908933
transform 1 0 20640 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1354
timestamp 1626908933
transform 1 0 20976 0 1 16761
box -32 -32 32 32
use M1M2_PR  M1M2_PR_586
timestamp 1626908933
transform 1 0 20976 0 1 16761
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_814
timestamp 1626908933
transform 1 0 21504 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_245
timestamp 1626908933
transform 1 0 21504 0 -1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_206
timestamp 1626908933
transform 1 0 21936 0 1 16539
box -32 -32 32 32
use M1M2_PR  M1M2_PR_974
timestamp 1626908933
transform 1 0 21936 0 1 16539
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_75
timestamp 1626908933
transform 1 0 21888 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_705
timestamp 1626908933
transform 1 0 21888 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_205
timestamp 1626908933
transform 1 0 21936 0 1 16909
box -32 -32 32 32
use M1M2_PR  M1M2_PR_973
timestamp 1626908933
transform 1 0 21936 0 1 16909
box -32 -32 32 32
use L1M1_PR  L1M1_PR_253
timestamp 1626908933
transform 1 0 22128 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1041
timestamp 1626908933
transform 1 0 22128 0 1 16539
box -29 -23 29 23
use L1M1_PR  L1M1_PR_652
timestamp 1626908933
transform 1 0 22224 0 1 16983
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1440
timestamp 1626908933
transform 1 0 22224 0 1 16983
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_5
timestamp 1626908933
transform 1 0 21984 0 -1 17316
box -38 -49 518 715
use sky130_fd_sc_hs__einvp_1  sky130_fd_sc_hs__einvp_1_15
timestamp 1626908933
transform 1 0 21984 0 -1 17316
box -38 -49 518 715
use L1M1_PR  L1M1_PR_1039
timestamp 1626908933
transform 1 0 22608 0 1 16835
box -29 -23 29 23
use L1M1_PR  L1M1_PR_251
timestamp 1626908933
transform 1 0 22608 0 1 16835
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_816
timestamp 1626908933
transform 1 0 22656 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_246
timestamp 1626908933
transform 1 0 22656 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_704
timestamp 1626908933
transform 1 0 22560 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_74
timestamp 1626908933
transform 1 0 22560 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_307
timestamp 1626908933
transform 1 0 22464 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_48
timestamp 1626908933
transform 1 0 22464 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_782
timestamp 1626908933
transform 1 0 23424 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_213
timestamp 1626908933
transform 1 0 23424 0 -1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1362
timestamp 1626908933
transform 1 0 24336 0 1 17131
box -32 -32 32 32
use M1M2_PR  M1M2_PR_594
timestamp 1626908933
transform 1 0 24336 0 1 17131
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_703
timestamp 1626908933
transform 1 0 23808 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_73
timestamp 1626908933
transform 1 0 23808 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_795
timestamp 1626908933
transform 1 0 23904 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_225
timestamp 1626908933
transform 1 0 23904 0 -1 17316
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_323
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_35
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_302
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_32
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_302
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_32
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_302
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_32
timestamp 1626908933
transform 1 0 24600 0 1 16650
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_420
timestamp 1626908933
transform 1 0 24672 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_52
timestamp 1626908933
transform 1 0 24672 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_199
timestamp 1626908933
transform 1 0 24864 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_768
timestamp 1626908933
transform 1 0 24864 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_774
timestamp 1626908933
transform 1 0 25248 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_204
timestamp 1626908933
transform 1 0 25248 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_746
timestamp 1626908933
transform 1 0 26016 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_177
timestamp 1626908933
transform 1 0 26016 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_702
timestamp 1626908933
transform 1 0 26400 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_72
timestamp 1626908933
transform 1 0 26400 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_752
timestamp 1626908933
transform 1 0 26496 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_182
timestamp 1626908933
transform 1 0 26496 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_51
timestamp 1626908933
transform 1 0 27552 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_419
timestamp 1626908933
transform 1 0 27552 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_47
timestamp 1626908933
transform 1 0 27456 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_306
timestamp 1626908933
transform 1 0 27456 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_71
timestamp 1626908933
transform 1 0 27264 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_587
timestamp 1626908933
transform 1 0 27360 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_701
timestamp 1626908933
transform 1 0 27264 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1217
timestamp 1626908933
transform 1 0 27360 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_70
timestamp 1626908933
transform 1 0 27744 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_700
timestamp 1626908933
transform 1 0 27744 0 -1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_602
timestamp 1626908933
transform 1 0 27696 0 1 16983
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1370
timestamp 1626908933
transform 1 0 27696 0 1 16983
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_158
timestamp 1626908933
transform 1 0 27840 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_728
timestamp 1626908933
transform 1 0 27840 0 -1 17316
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_307
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_19
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_17
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_287
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_17
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_287
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_17
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_287
timestamp 1626908933
transform 1 0 28600 0 1 16650
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_140
timestamp 1626908933
transform 1 0 28608 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_709
timestamp 1626908933
transform 1 0 28608 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_699
timestamp 1626908933
transform 1 0 28992 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_69
timestamp 1626908933
transform 1 0 28992 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_704
timestamp 1626908933
transform 1 0 29088 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_134
timestamp 1626908933
transform 1 0 29088 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_698
timestamp 1626908933
transform 1 0 29856 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_68
timestamp 1626908933
transform 1 0 29856 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_688
timestamp 1626908933
transform 1 0 29952 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_119
timestamp 1626908933
transform 1 0 29952 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_679
timestamp 1626908933
transform 1 0 30336 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_109
timestamp 1626908933
transform 1 0 30336 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_418
timestamp 1626908933
transform 1 0 31104 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_50
timestamp 1626908933
transform 1 0 31104 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_657
timestamp 1626908933
transform 1 0 31296 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_88
timestamp 1626908933
transform 1 0 31296 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_649
timestamp 1626908933
transform 1 0 31680 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_79
timestamp 1626908933
transform 1 0 31680 0 -1 17316
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_291
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_3
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_272
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_2
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_272
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_2
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_272
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_2
timestamp 1626908933
transform 1 0 32600 0 1 16650
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_305
timestamp 1626908933
transform 1 0 32448 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_46
timestamp 1626908933
transform 1 0 32448 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_55
timestamp 1626908933
transform 1 0 32544 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_624
timestamp 1626908933
transform 1 0 32544 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_619
timestamp 1626908933
transform 1 0 32928 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_49
timestamp 1626908933
transform 1 0 32928 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_697
timestamp 1626908933
transform 1 0 33696 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_67
timestamp 1626908933
transform 1 0 33696 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_591
timestamp 1626908933
transform 1 0 33792 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_22
timestamp 1626908933
transform 1 0 33792 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_589
timestamp 1626908933
transform 1 0 34176 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_19
timestamp 1626908933
transform 1 0 34176 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_2
timestamp 1626908933
transform 1 0 34944 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_572
timestamp 1626908933
transform 1 0 34944 0 -1 17316
box -38 -49 806 715
use M2M3_PR  M2M3_PR_101
timestamp 1626908933
transform 1 0 48 0 1 17849
box -33 -37 33 37
use M2M3_PR  M2M3_PR_42
timestamp 1626908933
transform 1 0 48 0 1 17849
box -33 -37 33 37
use M1M2_PR  M1M2_PR_1405
timestamp 1626908933
transform 1 0 48 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_637
timestamp 1626908933
transform 1 0 48 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_45
timestamp 1626908933
transform 1 0 288 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_304
timestamp 1626908933
transform 1 0 288 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_66
timestamp 1626908933
transform 1 0 384 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_696
timestamp 1626908933
transform 1 0 384 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_65
timestamp 1626908933
transform 1 0 864 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_695
timestamp 1626908933
transform 1 0 864 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_565
timestamp 1626908933
transform 1 0 480 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1134
timestamp 1626908933
transform 1 0 480 0 1 17316
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_130
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_418
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_588
timestamp 1626908933
transform 1 0 960 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1218
timestamp 1626908933
transform 1 0 960 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_165
timestamp 1626908933
transform 1 0 1104 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_933
timestamp 1626908933
transform 1 0 1104 0 1 17871
box -32 -32 32 32
use L1M1_PR  L1M1_PR_207
timestamp 1626908933
transform 1 0 1200 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_212
timestamp 1626908933
transform 1 0 1008 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_995
timestamp 1626908933
transform 1 0 1200 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1000
timestamp 1626908933
transform 1 0 1008 0 1 17871
box -29 -23 29 23
use M1M2_PR  M1M2_PR_161
timestamp 1626908933
transform 1 0 1296 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_929
timestamp 1626908933
transform 1 0 1296 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_160
timestamp 1626908933
transform 1 0 1296 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_928
timestamp 1626908933
transform 1 0 1296 0 1 17723
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_0
timestamp 1626908933
transform 1 0 1056 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_10
timestamp 1626908933
transform 1 0 1056 0 1 17316
box -38 -49 710 715
use L1M1_PR  L1M1_PR_204
timestamp 1626908933
transform 1 0 1488 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_633
timestamp 1626908933
transform 1 0 1584 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_992
timestamp 1626908933
transform 1 0 1488 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1421
timestamp 1626908933
transform 1 0 1584 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_549
timestamp 1626908933
transform 1 0 1728 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1118
timestamp 1626908933
transform 1 0 1728 0 1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_562
timestamp 1626908933
transform 1 0 2352 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1330
timestamp 1626908933
transform 1 0 2352 0 1 17427
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_553
timestamp 1626908933
transform 1 0 2112 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1123
timestamp 1626908933
transform 1 0 2112 0 1 17316
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_257
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_527
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_257
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_527
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_257
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_527
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_562
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_274
timestamp 1626908933
transform 1 0 2600 0 1 17316
box -200 -142 200 178
use M1M2_PR  M1M2_PR_170
timestamp 1626908933
transform 1 0 2928 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_938
timestamp 1626908933
transform 1 0 2928 0 1 17871
box -32 -32 32 32
use L1M1_PR  L1M1_PR_217
timestamp 1626908933
transform 1 0 2832 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1005
timestamp 1626908933
transform 1 0 2832 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_203
timestamp 1626908933
transform 1 0 3024 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_991
timestamp 1626908933
transform 1 0 3024 0 1 17723
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_1
timestamp 1626908933
transform 1 0 2880 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_11
timestamp 1626908933
transform 1 0 2880 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_528
timestamp 1626908933
transform 1 0 3552 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1097
timestamp 1626908933
transform 1 0 3552 0 1 17316
box -38 -49 422 715
use L1M1_PR  L1M1_PR_199
timestamp 1626908933
transform 1 0 3312 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_637
timestamp 1626908933
transform 1 0 3408 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_987
timestamp 1626908933
transform 1 0 3312 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1425
timestamp 1626908933
transform 1 0 3408 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_739
timestamp 1626908933
transform 1 0 4080 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1527
timestamp 1626908933
transform 1 0 4080 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_712
timestamp 1626908933
transform 1 0 3792 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1480
timestamp 1626908933
transform 1 0 3792 0 1 17649
box -32 -32 32 32
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_52
timestamp 1626908933
transform 1 0 3936 0 1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_132
timestamp 1626908933
transform 1 0 3936 0 1 17316
box -38 -49 902 715
use M1M2_PR  M1M2_PR_1341
timestamp 1626908933
transform 1 0 4464 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_573
timestamp 1626908933
transform 1 0 4464 0 1 17427
box -32 -32 32 32
use L1M1_PR  L1M1_PR_964
timestamp 1626908933
transform 1 0 4464 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_176
timestamp 1626908933
transform 1 0 4464 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_908
timestamp 1626908933
transform 1 0 4272 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_140
timestamp 1626908933
transform 1 0 4272 0 1 17649
box -32 -32 32 32
use M2M3_PR  M2M3_PR_91
timestamp 1626908933
transform 1 0 4464 0 1 17483
box -33 -37 33 37
use M2M3_PR  M2M3_PR_32
timestamp 1626908933
transform 1 0 4464 0 1 17483
box -33 -37 33 37
use osc_core_VIA4  osc_core_VIA4_402
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_114
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_351
timestamp 1626908933
transform 1 0 4800 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_719
timestamp 1626908933
transform 1 0 4800 0 1 17316
box -38 -49 230 715
use M1M2_PR  M1M2_PR_754
timestamp 1626908933
transform 1 0 4848 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1522
timestamp 1626908933
transform 1 0 4848 0 1 17205
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_44
timestamp 1626908933
transform 1 0 4992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_303
timestamp 1626908933
transform 1 0 4992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_352
timestamp 1626908933
transform 1 0 5472 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_720
timestamp 1626908933
transform 1 0 5472 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_589
timestamp 1626908933
transform 1 0 5664 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1219
timestamp 1626908933
transform 1 0 5664 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_233
timestamp 1626908933
transform 1 0 5808 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1001
timestamp 1626908933
transform 1 0 5808 0 1 17871
box -32 -32 32 32
use L1M1_PR  L1M1_PR_288
timestamp 1626908933
transform 1 0 5712 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1076
timestamp 1626908933
transform 1 0 5712 0 1 17871
box -29 -23 29 23
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_7
timestamp 1626908933
transform 1 0 5088 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_16
timestamp 1626908933
transform 1 0 5088 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_8
timestamp 1626908933
transform 1 0 5760 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_18
timestamp 1626908933
transform 1 0 5760 0 1 17316
box -38 -49 710 715
use M1M2_PR  M1M2_PR_997
timestamp 1626908933
transform 1 0 6000 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_229
timestamp 1626908933
transform 1 0 6000 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1068
timestamp 1626908933
transform 1 0 6192 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_280
timestamp 1626908933
transform 1 0 6192 0 1 17205
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1398
timestamp 1626908933
transform 1 0 6192 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_630
timestamp 1626908933
transform 1 0 6192 0 1 17427
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1071
timestamp 1626908933
transform 1 0 5904 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_283
timestamp 1626908933
transform 1 0 5904 0 1 17723
box -29 -23 29 23
use M1M2_PR  M1M2_PR_996
timestamp 1626908933
transform 1 0 6000 0 1 17723
box -32 -32 32 32
use M1M2_PR  M1M2_PR_228
timestamp 1626908933
transform 1 0 6000 0 1 17723
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_242
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_512
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_242
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_512
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_242
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_512
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -49 200 49
use L1M1_PR  L1M1_PR_665
timestamp 1626908933
transform 1 0 6288 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1453
timestamp 1626908933
transform 1 0 6288 0 1 17427
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_258
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_546
timestamp 1626908933
transform 1 0 6600 0 1 17316
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_417
timestamp 1626908933
transform 1 0 6432 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_49
timestamp 1626908933
transform 1 0 6432 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_504
timestamp 1626908933
transform 1 0 6624 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1074
timestamp 1626908933
transform 1 0 6624 0 1 17316
box -38 -49 806 715
use M2M3_PR  M2M3_PR_100
timestamp 1626908933
transform 1 0 6864 0 1 17727
box -33 -37 33 37
use M2M3_PR  M2M3_PR_41
timestamp 1626908933
transform 1 0 6864 0 1 17727
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_48
timestamp 1626908933
transform 1 0 7392 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_416
timestamp 1626908933
transform 1 0 7392 0 1 17316
box -38 -49 230 715
use L1M1_PR  L1M1_PR_279
timestamp 1626908933
transform 1 0 7728 0 1 17723
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1067
timestamp 1626908933
transform 1 0 7728 0 1 17723
box -29 -23 29 23
use M1M2_PR  M1M2_PR_237
timestamp 1626908933
transform 1 0 7632 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1005
timestamp 1626908933
transform 1 0 7632 0 1 17871
box -32 -32 32 32
use L1M1_PR  L1M1_PR_293
timestamp 1626908933
transform 1 0 7536 0 1 17871
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1081
timestamp 1626908933
transform 1 0 7536 0 1 17871
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_9
timestamp 1626908933
transform 1 0 7584 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_19
timestamp 1626908933
transform 1 0 7584 0 1 17316
box -38 -49 710 715
use osc_core_VIA4  osc_core_VIA4_386
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_98
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -142 200 178
use L1M1_PR  L1M1_PR_1063
timestamp 1626908933
transform 1 0 8016 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_275
timestamp 1626908933
transform 1 0 8016 0 1 17205
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1058
timestamp 1626908933
transform 1 0 8256 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_488
timestamp 1626908933
transform 1 0 8256 0 1 17316
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1457
timestamp 1626908933
transform 1 0 8112 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_669
timestamp 1626908933
transform 1 0 8112 0 1 17427
box -29 -23 29 23
use M1M2_PR  M1M2_PR_77
timestamp 1626908933
transform 1 0 9648 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_845
timestamp 1626908933
transform 1 0 9648 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_89
timestamp 1626908933
transform 1 0 9648 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_877
timestamp 1626908933
transform 1 0 9648 0 1 17649
box -29 -23 29 23
use M1M2_PR  M1M2_PR_717
timestamp 1626908933
transform 1 0 9264 0 1 17649
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1485
timestamp 1626908933
transform 1 0 9264 0 1 17649
box -32 -32 32 32
use L1M1_PR  L1M1_PR_748
timestamp 1626908933
transform 1 0 9264 0 1 17649
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1536
timestamp 1626908933
transform 1 0 9264 0 1 17649
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_42
timestamp 1626908933
transform 1 0 9024 0 1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_122
timestamp 1626908933
transform 1 0 9024 0 1 17316
box -38 -49 902 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_43
timestamp 1626908933
transform 1 0 9984 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_302
timestamp 1626908933
transform 1 0 9984 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_590
timestamp 1626908933
transform 1 0 9888 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1220
timestamp 1626908933
transform 1 0 9888 0 1 17316
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_530
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_242
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_227
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_497
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_227
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_497
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_227
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_497
timestamp 1626908933
transform 1 0 10600 0 1 17316
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_459
timestamp 1626908933
transform 1 0 10464 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1029
timestamp 1626908933
transform 1 0 10464 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_444
timestamp 1626908933
transform 1 0 10080 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1013
timestamp 1626908933
transform 1 0 10080 0 1 17316
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1018
timestamp 1626908933
transform 1 0 11376 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_230
timestamp 1626908933
transform 1 0 11376 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_12
timestamp 1626908933
transform 1 0 11328 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_2
timestamp 1626908933
transform 1 0 11328 0 1 17316
box -38 -49 710 715
use M1M2_PR  M1M2_PR_950
timestamp 1626908933
transform 1 0 11376 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_182
timestamp 1626908933
transform 1 0 11376 0 1 17575
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1221
timestamp 1626908933
transform 1 0 11232 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_591
timestamp 1626908933
transform 1 0 11232 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_641
timestamp 1626908933
transform 1 0 11856 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1429
timestamp 1626908933
transform 1 0 11856 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_223
timestamp 1626908933
transform 1 0 11760 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1011
timestamp 1626908933
transform 1 0 11760 0 1 17205
box -29 -23 29 23
use M1M2_PR  M1M2_PR_178
timestamp 1626908933
transform 1 0 11664 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_946
timestamp 1626908933
transform 1 0 11664 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_177
timestamp 1626908933
transform 1 0 11664 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_945
timestamp 1626908933
transform 1 0 11664 0 1 17797
box -32 -32 32 32
use L1M1_PR  L1M1_PR_226
timestamp 1626908933
transform 1 0 11472 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1014
timestamp 1626908933
transform 1 0 11472 0 1 17797
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_414
timestamp 1626908933
transform 1 0 12000 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_983
timestamp 1626908933
transform 1 0 12000 0 1 17316
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_370
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_82
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1008
timestamp 1626908933
transform 1 0 12384 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_438
timestamp 1626908933
transform 1 0 12384 0 1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_187
timestamp 1626908933
transform 1 0 13104 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_955
timestamp 1626908933
transform 1 0 13104 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_186
timestamp 1626908933
transform 1 0 13104 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_954
timestamp 1626908933
transform 1 0 13104 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_222
timestamp 1626908933
transform 1 0 13296 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1010
timestamp 1626908933
transform 1 0 13296 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_236
timestamp 1626908933
transform 1 0 13200 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1024
timestamp 1626908933
transform 1 0 13200 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_3
timestamp 1626908933
transform 1 0 13152 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_13
timestamp 1626908933
transform 1 0 13152 0 1 17316
box -38 -49 710 715
use L1M1_PR  L1M1_PR_232
timestamp 1626908933
transform 1 0 13680 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_645
timestamp 1626908933
transform 1 0 13680 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1020
timestamp 1626908933
transform 1 0 13680 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1433
timestamp 1626908933
transform 1 0 13680 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_218
timestamp 1626908933
transform 1 0 13584 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1006
timestamp 1626908933
transform 1 0 13584 0 1 17131
box -29 -23 29 23
use M1M2_PR  M1M2_PR_588
timestamp 1626908933
transform 1 0 13872 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1356
timestamp 1626908933
transform 1 0 13872 0 1 17427
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_372
timestamp 1626908933
transform 1 0 13824 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_941
timestamp 1626908933
transform 1 0 13824 0 1 17316
box -38 -49 422 715
use osc_core_VIA5  osc_core_VIA5_212
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_482
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_212
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_482
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_212
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_482
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -49 200 49
use M1M2_PR  M1M2_PR_582
timestamp 1626908933
transform 1 0 14352 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1350
timestamp 1626908933
transform 1 0 14352 0 1 17427
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_514
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_226
timestamp 1626908933
transform 1 0 14600 0 1 17316
box -200 -142 200 178
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_42
timestamp 1626908933
transform 1 0 14976 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_301
timestamp 1626908933
transform 1 0 14976 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_410
timestamp 1626908933
transform 1 0 14208 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_980
timestamp 1626908933
transform 1 0 14208 0 1 17316
box -38 -49 806 715
use M2M3_PR  M2M3_PR_90
timestamp 1626908933
transform 1 0 15024 0 1 17483
box -33 -37 33 37
use M2M3_PR  M2M3_PR_31
timestamp 1626908933
transform 1 0 15024 0 1 17483
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_415
timestamp 1626908933
transform 1 0 15072 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_47
timestamp 1626908933
transform 1 0 15072 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_953
timestamp 1626908933
transform 1 0 15264 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_383
timestamp 1626908933
transform 1 0 15264 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_16
timestamp 1626908933
transform 1 0 16032 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_6
timestamp 1626908933
transform 1 0 16032 0 1 17316
box -38 -49 710 715
use M1M2_PR  M1M2_PR_985
timestamp 1626908933
transform 1 0 16272 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_217
timestamp 1626908933
transform 1 0 16272 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1050
timestamp 1626908933
transform 1 0 16464 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_262
timestamp 1626908933
transform 1 0 16464 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1056
timestamp 1626908933
transform 1 0 16080 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_268
timestamp 1626908933
transform 1 0 16080 0 1 17575
box -29 -23 29 23
use M1M2_PR  M1M2_PR_984
timestamp 1626908933
transform 1 0 16272 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_216
timestamp 1626908933
transform 1 0 16272 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1052
timestamp 1626908933
transform 1 0 16176 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_264
timestamp 1626908933
transform 1 0 16176 0 1 17797
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_66
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_354
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -142 200 178
use M1M2_PR  M1M2_PR_980
timestamp 1626908933
transform 1 0 16464 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_212
timestamp 1626908933
transform 1 0 16464 0 1 17797
box -32 -32 32 32
use L1M1_PR  L1M1_PR_265
timestamp 1626908933
transform 1 0 16560 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_657
timestamp 1626908933
transform 1 0 16560 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1053
timestamp 1626908933
transform 1 0 16560 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1445
timestamp 1626908933
transform 1 0 16560 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_46
timestamp 1626908933
transform 1 0 16704 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_414
timestamp 1626908933
transform 1 0 16704 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_356
timestamp 1626908933
transform 1 0 16896 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_926
timestamp 1626908933
transform 1 0 16896 0 1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_976
timestamp 1626908933
transform 1 0 17616 0 1 17871
box -32 -32 32 32
use M1M2_PR  M1M2_PR_208
timestamp 1626908933
transform 1 0 17616 0 1 17871
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_413
timestamp 1626908933
transform 1 0 17664 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_45
timestamp 1626908933
transform 1 0 17664 0 1 17316
box -38 -49 230 715
use L1M1_PR  L1M1_PR_1062
timestamp 1626908933
transform 1 0 17904 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_274
timestamp 1626908933
transform 1 0 17904 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_17
timestamp 1626908933
transform 1 0 17856 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_7
timestamp 1626908933
transform 1 0 17856 0 1 17316
box -38 -49 710 715
use M1M2_PR  M1M2_PR_990
timestamp 1626908933
transform 1 0 17808 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_222
timestamp 1626908933
transform 1 0 17808 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_661
timestamp 1626908933
transform 1 0 18384 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1449
timestamp 1626908933
transform 1 0 18384 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_256
timestamp 1626908933
transform 1 0 18288 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1044
timestamp 1626908933
transform 1 0 18288 0 1 17131
box -29 -23 29 23
use L1M1_PR  L1M1_PR_259
timestamp 1626908933
transform 1 0 18000 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1047
timestamp 1626908933
transform 1 0 18000 0 1 17797
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_210
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_498
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_467
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_197
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_467
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_197
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_467
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_197
timestamp 1626908933
transform 1 0 18600 0 1 17316
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_694
timestamp 1626908933
transform 1 0 18720 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_64
timestamp 1626908933
transform 1 0 18720 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_412
timestamp 1626908933
transform 1 0 18528 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_44
timestamp 1626908933
transform 1 0 18528 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_333
timestamp 1626908933
transform 1 0 18816 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_903
timestamp 1626908933
transform 1 0 18816 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_846
timestamp 1626908933
transform 1 0 19584 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_277
timestamp 1626908933
transform 1 0 19584 0 1 17316
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1378
timestamp 1626908933
transform 1 0 18864 0 1 17501
box -32 -32 32 32
use M1M2_PR  M1M2_PR_610
timestamp 1626908933
transform 1 0 18864 0 1 17501
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_592
timestamp 1626908933
transform 1 0 20064 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1222
timestamp 1626908933
transform 1 0 20064 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_41
timestamp 1626908933
transform 1 0 19968 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_300
timestamp 1626908933
transform 1 0 19968 0 1 17316
box -38 -49 134 715
use M1M2_PR  M1M2_PR_621
timestamp 1626908933
transform 1 0 19920 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1389
timestamp 1626908933
transform 1 0 19920 0 1 17427
box -32 -32 32 32
use M2M3_PR  M2M3_PR_36
timestamp 1626908933
transform 1 0 19920 0 1 17483
box -33 -37 33 37
use M2M3_PR  M2M3_PR_95
timestamp 1626908933
transform 1 0 19920 0 1 17483
box -33 -37 33 37
use M1M2_PR  M1M2_PR_197
timestamp 1626908933
transform 1 0 20400 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_965
timestamp 1626908933
transform 1 0 20400 0 1 17575
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_338
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_50
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -142 200 178
use L1M1_PR  L1M1_PR_245
timestamp 1626908933
transform 1 0 20304 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_249
timestamp 1626908933
transform 1 0 20208 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1033
timestamp 1626908933
transform 1 0 20304 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1037
timestamp 1626908933
transform 1 0 20208 0 1 17575
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_4
timestamp 1626908933
transform 1 0 20160 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_14
timestamp 1626908933
transform 1 0 20160 0 1 17316
box -38 -49 710 715
use M1M2_PR  M1M2_PR_960
timestamp 1626908933
transform 1 0 20592 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_192
timestamp 1626908933
transform 1 0 20592 0 1 17797
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1437
timestamp 1626908933
transform 1 0 20688 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1030
timestamp 1626908933
transform 1 0 20592 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_649
timestamp 1626908933
transform 1 0 20688 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_242
timestamp 1626908933
transform 1 0 20592 0 1 17205
box -29 -23 29 23
use M1M2_PR  M1M2_PR_961
timestamp 1626908933
transform 1 0 20592 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_193
timestamp 1626908933
transform 1 0 20592 0 1 17205
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_818
timestamp 1626908933
transform 1 0 20832 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_249
timestamp 1626908933
transform 1 0 20832 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_843
timestamp 1626908933
transform 1 0 21216 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_273
timestamp 1626908933
transform 1 0 21216 0 1 17316
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1364
timestamp 1626908933
transform 1 0 21744 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_596
timestamp 1626908933
transform 1 0 21744 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_958
timestamp 1626908933
transform 1 0 22320 0 1 17205
box -32 -32 32 32
use M1M2_PR  M1M2_PR_190
timestamp 1626908933
transform 1 0 22320 0 1 17205
box -32 -32 32 32
use L1M1_PR  L1M1_PR_237
timestamp 1626908933
transform 1 0 22416 0 1 17205
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1025
timestamp 1626908933
transform 1 0 22416 0 1 17205
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_182
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_452
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_182
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_452
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_182
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_452
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_194
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_482
timestamp 1626908933
transform 1 0 22600 0 1 17316
box -200 -142 200 178
use M1M2_PR  M1M2_PR_204
timestamp 1626908933
transform 1 0 21936 0 1 17575
box -32 -32 32 32
use M1M2_PR  M1M2_PR_972
timestamp 1626908933
transform 1 0 21936 0 1 17575
box -32 -32 32 32
use L1M1_PR  L1M1_PR_240
timestamp 1626908933
transform 1 0 22128 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_255
timestamp 1626908933
transform 1 0 22032 0 1 17575
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1028
timestamp 1626908933
transform 1 0 22128 0 1 17797
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1043
timestamp 1626908933
transform 1 0 22032 0 1 17575
box -29 -23 29 23
use M1M2_PR  M1M2_PR_189
timestamp 1626908933
transform 1 0 22320 0 1 17797
box -32 -32 32 32
use M1M2_PR  M1M2_PR_957
timestamp 1626908933
transform 1 0 22320 0 1 17797
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_5
timestamp 1626908933
transform 1 0 21984 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__einvp_2  sky130_fd_sc_hs__einvp_2_15
timestamp 1626908933
transform 1 0 21984 0 1 17316
box -38 -49 710 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_801
timestamp 1626908933
transform 1 0 22944 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_232
timestamp 1626908933
transform 1 0 22944 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_411
timestamp 1626908933
transform 1 0 22752 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_43
timestamp 1626908933
transform 1 0 22752 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_299
timestamp 1626908933
transform 1 0 22656 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_40
timestamp 1626908933
transform 1 0 22656 0 1 17316
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1441
timestamp 1626908933
transform 1 0 22512 0 1 17427
box -29 -23 29 23
use L1M1_PR  L1M1_PR_653
timestamp 1626908933
transform 1 0 22512 0 1 17427
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_813
timestamp 1626908933
transform 1 0 23328 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_243
timestamp 1626908933
transform 1 0 23328 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_693
timestamp 1626908933
transform 1 0 24096 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_63
timestamp 1626908933
transform 1 0 24096 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_792
timestamp 1626908933
transform 1 0 24192 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_222
timestamp 1626908933
transform 1 0 24192 0 1 17316
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_322
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_34
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_410
timestamp 1626908933
transform 1 0 25056 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_42
timestamp 1626908933
transform 1 0 25056 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_298
timestamp 1626908933
transform 1 0 24960 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_39
timestamp 1626908933
transform 1 0 24960 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_773
timestamp 1626908933
transform 1 0 25248 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_203
timestamp 1626908933
transform 1 0 25248 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_745
timestamp 1626908933
transform 1 0 26016 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_176
timestamp 1626908933
transform 1 0 26016 0 1 17316
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_466
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_178
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_437
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_167
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_437
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_167
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_437
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_167
timestamp 1626908933
transform 1 0 26600 0 1 17316
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_692
timestamp 1626908933
transform 1 0 26400 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_62
timestamp 1626908933
transform 1 0 26400 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_181
timestamp 1626908933
transform 1 0 26496 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_751
timestamp 1626908933
transform 1 0 26496 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_727
timestamp 1626908933
transform 1 0 27840 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_157
timestamp 1626908933
transform 1 0 27840 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_409
timestamp 1626908933
transform 1 0 27264 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_41
timestamp 1626908933
transform 1 0 27264 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_731
timestamp 1626908933
transform 1 0 27456 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_162
timestamp 1626908933
transform 1 0 27456 0 1 17316
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_18
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_306
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -142 200 178
use M1M2_PR  M1M2_PR_1371
timestamp 1626908933
transform 1 0 28272 0 1 17427
box -32 -32 32 32
use M1M2_PR  M1M2_PR_603
timestamp 1626908933
transform 1 0 28272 0 1 17427
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_708
timestamp 1626908933
transform 1 0 28608 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_139
timestamp 1626908933
transform 1 0 28608 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_691
timestamp 1626908933
transform 1 0 28992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_61
timestamp 1626908933
transform 1 0 28992 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_703
timestamp 1626908933
transform 1 0 29088 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_133
timestamp 1626908933
transform 1 0 29088 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1223
timestamp 1626908933
transform 1 0 29856 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_593
timestamp 1626908933
transform 1 0 29856 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_60
timestamp 1626908933
transform 1 0 30240 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_690
timestamp 1626908933
transform 1 0 30240 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_38
timestamp 1626908933
transform 1 0 29952 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_297
timestamp 1626908933
transform 1 0 29952 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_40
timestamp 1626908933
transform 1 0 30048 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_408
timestamp 1626908933
transform 1 0 30048 0 1 17316
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_152
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_422
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_152
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_422
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_152
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_422
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_162
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_450
timestamp 1626908933
transform 1 0 30600 0 1 17316
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_108
timestamp 1626908933
transform 1 0 30336 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_678
timestamp 1626908933
transform 1 0 30336 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_407
timestamp 1626908933
transform 1 0 31104 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_39
timestamp 1626908933
transform 1 0 31104 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_656
timestamp 1626908933
transform 1 0 31296 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_87
timestamp 1626908933
transform 1 0 31296 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_648
timestamp 1626908933
transform 1 0 31680 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_78
timestamp 1626908933
transform 1 0 31680 0 1 17316
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_290
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_2
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_689
timestamp 1626908933
transform 1 0 32448 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_59
timestamp 1626908933
transform 1 0 32448 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_623
timestamp 1626908933
transform 1 0 32544 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_54
timestamp 1626908933
transform 1 0 32544 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_618
timestamp 1626908933
transform 1 0 32928 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_48
timestamp 1626908933
transform 1 0 32928 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_688
timestamp 1626908933
transform 1 0 33696 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_58
timestamp 1626908933
transform 1 0 33696 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_590
timestamp 1626908933
transform 1 0 33792 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_21
timestamp 1626908933
transform 1 0 33792 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_588
timestamp 1626908933
transform 1 0 34176 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_18
timestamp 1626908933
transform 1 0 34176 0 1 17316
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_407
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_137
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_407
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_137
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_407
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_137
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_146
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_434
timestamp 1626908933
transform 1 0 34600 0 1 17316
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_571
timestamp 1626908933
transform 1 0 35040 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_2
timestamp 1626908933
transform 1 0 35040 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_296
timestamp 1626908933
transform 1 0 34944 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_37
timestamp 1626908933
transform 1 0 34944 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_721
timestamp 1626908933
transform 1 0 35424 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_353
timestamp 1626908933
transform 1 0 35424 0 1 17316
box -38 -49 230 715
use M2M3_PR  M2M3_PR_94
timestamp 1626908933
transform 1 0 35184 0 1 17239
box -33 -37 33 37
use M2M3_PR  M2M3_PR_35
timestamp 1626908933
transform 1 0 35184 0 1 17239
box -33 -37 33 37
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1224
timestamp 1626908933
transform 1 0 35616 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_594
timestamp 1626908933
transform 1 0 35616 0 1 17316
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_391
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_121
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_391
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_121
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_391
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_121
timestamp 1626908933
transform 1 0 600 0 1 17982
box -200 -49 200 49
use M1M2_PR  M1M2_PR_1403
timestamp 1626908933
transform 1 0 48 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_635
timestamp 1626908933
transform 1 0 48 0 1 18537
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_678
timestamp 1626908933
transform 1 0 384 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_48
timestamp 1626908933
transform 1 0 384 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_288
timestamp 1626908933
transform 1 0 288 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_29
timestamp 1626908933
transform 1 0 288 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1133
timestamp 1626908933
transform 1 0 480 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_564
timestamp 1626908933
transform 1 0 480 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_677
timestamp 1626908933
transform 1 0 864 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_47
timestamp 1626908933
transform 1 0 864 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1230
timestamp 1626908933
transform 1 0 960 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_600
timestamp 1626908933
transform 1 0 960 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_994
timestamp 1626908933
transform 1 0 1200 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_206
timestamp 1626908933
transform 1 0 1200 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_999
timestamp 1626908933
transform 1 0 1104 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_211
timestamp 1626908933
transform 1 0 1104 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_932
timestamp 1626908933
transform 1 0 1104 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_164
timestamp 1626908933
transform 1 0 1104 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_927
timestamp 1626908933
transform 1 0 1296 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_159
timestamp 1626908933
transform 1 0 1296 0 1 18167
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_567
timestamp 1626908933
transform 1 0 288 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1137
timestamp 1626908933
transform 1 0 288 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_0
timestamp 1626908933
transform 1 0 1056 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_10
timestamp 1626908933
transform 1 0 1056 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_10
timestamp 1626908933
transform 1 0 1056 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_0
timestamp 1626908933
transform 1 0 1056 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_354
timestamp 1626908933
transform 1 0 2208 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_722
timestamp 1626908933
transform 1 0 2208 0 -1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_634
timestamp 1626908933
transform 1 0 2160 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1422
timestamp 1626908933
transform 1 0 2160 0 1 18389
box -29 -23 29 23
use osc_core_VIA7  osc_core_VIA7_526
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_256
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_526
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_256
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_526
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_256
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_273
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_561
timestamp 1626908933
transform 1 0 2600 0 1 18648
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1225
timestamp 1626908933
transform 1 0 2400 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_595
timestamp 1626908933
transform 1 0 2400 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_295
timestamp 1626908933
transform 1 0 2496 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_36
timestamp 1626908933
transform 1 0 2496 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_723
timestamp 1626908933
transform 1 0 2592 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_355
timestamp 1626908933
transform 1 0 2592 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_596
timestamp 1626908933
transform 1 0 2784 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1226
timestamp 1626908933
transform 1 0 2784 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_202
timestamp 1626908933
transform 1 0 3024 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_990
timestamp 1626908933
transform 1 0 3024 0 1 18167
box -29 -23 29 23
use M1M2_PR  M1M2_PR_169
timestamp 1626908933
transform 1 0 2928 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_937
timestamp 1626908933
transform 1 0 2928 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_216
timestamp 1626908933
transform 1 0 2928 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1004
timestamp 1626908933
transform 1 0 2928 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_567
timestamp 1626908933
transform 1 0 3312 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1335
timestamp 1626908933
transform 1 0 3312 0 1 18389
box -32 -32 32 32
use M2M3_PR  M2M3_PR_34
timestamp 1626908933
transform 1 0 4176 0 1 18337
box -33 -37 33 37
use M2M3_PR  M2M3_PR_93
timestamp 1626908933
transform 1 0 4176 0 1 18337
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_356
timestamp 1626908933
transform 1 0 4032 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_724
timestamp 1626908933
transform 1 0 4032 0 -1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_638
timestamp 1626908933
transform 1 0 3984 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1426
timestamp 1626908933
transform 1 0 3984 0 1 18389
box -29 -23 29 23
use M1M2_PR  M1M2_PR_574
timestamp 1626908933
transform 1 0 4176 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1342
timestamp 1626908933
transform 1 0 4176 0 1 18389
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_1
timestamp 1626908933
transform 1 0 2880 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_11
timestamp 1626908933
transform 1 0 2880 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_11
timestamp 1626908933
transform 1 0 2880 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_1
timestamp 1626908933
transform 1 0 2880 0 1 18648
box -38 -49 1862 715
use osc_core_VIA7  osc_core_VIA7_376
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_106
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_376
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_106
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_376
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_106
timestamp 1626908933
transform 1 0 4600 0 1 17982
box -200 -49 200 49
use M1M2_PR  M1M2_PR_138
timestamp 1626908933
transform 1 0 4368 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_906
timestamp 1626908933
transform 1 0 4368 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_175
timestamp 1626908933
transform 1 0 4464 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_963
timestamp 1626908933
transform 1 0 4464 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_632
timestamp 1626908933
transform 1 0 4560 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1400
timestamp 1626908933
transform 1 0 4560 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_753
timestamp 1626908933
transform 1 0 4848 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1521
timestamp 1626908933
transform 1 0 4848 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_778
timestamp 1626908933
transform 1 0 4848 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1566
timestamp 1626908933
transform 1 0 4848 0 1 18315
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_728
timestamp 1626908933
transform 1 0 4704 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_360
timestamp 1626908933
transform 1 0 4704 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1227
timestamp 1626908933
transform 1 0 4224 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_597
timestamp 1626908933
transform 1 0 4224 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1231
timestamp 1626908933
transform 1 0 4896 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_601
timestamp 1626908933
transform 1 0 4896 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_287
timestamp 1626908933
transform 1 0 4992 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_28
timestamp 1626908933
transform 1 0 4992 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_406
timestamp 1626908933
transform 1 0 5184 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_38
timestamp 1626908933
transform 1 0 5184 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_729
timestamp 1626908933
transform 1 0 5472 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_361
timestamp 1626908933
transform 1 0 5472 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_17
timestamp 1626908933
transform 1 0 5088 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_8
timestamp 1626908933
transform 1 0 5088 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1079
timestamp 1626908933
transform 1 0 5376 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_510
timestamp 1626908933
transform 1 0 5376 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_63
timestamp 1626908933
transform -1 0 5184 0 -1 18648
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_143
timestamp 1626908933
transform -1 0 5184 0 -1 18648
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1232
timestamp 1626908933
transform 1 0 5664 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_602
timestamp 1626908933
transform 1 0 5664 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1074
timestamp 1626908933
transform 1 0 5808 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_286
timestamp 1626908933
transform 1 0 5808 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1000
timestamp 1626908933
transform 1 0 5808 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_232
timestamp 1626908933
transform 1 0 5808 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_995
timestamp 1626908933
transform 1 0 6000 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_227
timestamp 1626908933
transform 1 0 6000 0 1 18167
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1070
timestamp 1626908933
transform 1 0 6096 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_282
timestamp 1626908933
transform 1 0 6096 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_666
timestamp 1626908933
transform 1 0 6864 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1454
timestamp 1626908933
transform 1 0 6864 0 1 18389
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_241
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_511
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_241
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_511
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_241
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_511
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_545
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_257
timestamp 1626908933
transform 1 0 6600 0 1 18648
box -200 -142 200 178
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1061
timestamp 1626908933
transform 1 0 6912 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_492
timestamp 1626908933
transform 1 0 6912 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_8
timestamp 1626908933
transform 1 0 5760 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_18
timestamp 1626908933
transform 1 0 5760 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_18
timestamp 1626908933
transform 1 0 5760 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_8
timestamp 1626908933
transform 1 0 5760 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_357
timestamp 1626908933
transform 1 0 7296 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_725
timestamp 1626908933
transform 1 0 7296 0 -1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_236
timestamp 1626908933
transform 1 0 7632 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1004
timestamp 1626908933
transform 1 0 7632 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_35
timestamp 1626908933
transform 1 0 7488 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_294
timestamp 1626908933
transform 1 0 7488 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_634
timestamp 1626908933
transform 1 0 7440 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1402
timestamp 1626908933
transform 1 0 7440 0 1 18537
box -32 -32 32 32
use L1M1_PR  L1M1_PR_278
timestamp 1626908933
transform 1 0 7728 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1066
timestamp 1626908933
transform 1 0 7728 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_292
timestamp 1626908933
transform 1 0 7632 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1080
timestamp 1626908933
transform 1 0 7632 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_638
timestamp 1626908933
transform 1 0 8304 0 1 18389
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1406
timestamp 1626908933
transform 1 0 8304 0 1 18389
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_9
timestamp 1626908933
transform 1 0 7584 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_19
timestamp 1626908933
transform 1 0 7584 0 -1 18648
box -38 -49 1190 715
use osc_core_VIA7  osc_core_VIA7_361
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_91
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_361
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_91
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_361
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_91
timestamp 1626908933
transform 1 0 8600 0 1 17982
box -200 -49 200 49
use L1M1_PR  L1M1_PR_1458
timestamp 1626908933
transform 1 0 8688 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_670
timestamp 1626908933
transform 1 0 8688 0 1 18389
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1039
timestamp 1626908933
transform 1 0 8736 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_470
timestamp 1626908933
transform 1 0 8736 0 -1 18648
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1535
timestamp 1626908933
transform 1 0 9264 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_747
timestamp 1626908933
transform 1 0 9264 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1484
timestamp 1626908933
transform 1 0 9264 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_716
timestamp 1626908933
transform 1 0 9264 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_676
timestamp 1626908933
transform 1 0 9408 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_46
timestamp 1626908933
transform 1 0 9408 0 1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_876
timestamp 1626908933
transform 1 0 9648 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_88
timestamp 1626908933
transform 1 0 9648 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_844
timestamp 1626908933
transform 1 0 9648 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_76
timestamp 1626908933
transform 1 0 9648 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1031
timestamp 1626908933
transform 1 0 9504 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_462
timestamp 1626908933
transform 1 0 9504 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_40
timestamp 1626908933
transform 1 0 9120 0 -1 18648
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_120
timestamp 1626908933
transform 1 0 9120 0 -1 18648
box -38 -49 902 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_19
timestamp 1626908933
transform 1 0 7584 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_9
timestamp 1626908933
transform 1 0 7584 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_675
timestamp 1626908933
transform 1 0 9888 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_45
timestamp 1626908933
transform 1 0 9888 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_286
timestamp 1626908933
transform 1 0 9984 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_27
timestamp 1626908933
transform 1 0 9984 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_687
timestamp 1626908933
transform 1 0 9984 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_57
timestamp 1626908933
transform 1 0 9984 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1011
timestamp 1626908933
transform 1 0 10080 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_442
timestamp 1626908933
transform 1 0 10080 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1012
timestamp 1626908933
transform 1 0 10080 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_443
timestamp 1626908933
transform 1 0 10080 0 -1 18648
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_529
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_241
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_226
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_496
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_226
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_496
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_226
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_496
timestamp 1626908933
transform 1 0 10600 0 1 18648
box -200 -49 200 49
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_458
timestamp 1626908933
transform 1 0 10464 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1028
timestamp 1626908933
transform 1 0 10464 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_457
timestamp 1626908933
transform 1 0 10464 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1027
timestamp 1626908933
transform 1 0 10464 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1233
timestamp 1626908933
transform 1 0 11232 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_603
timestamp 1626908933
transform 1 0 11232 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_686
timestamp 1626908933
transform 1 0 11232 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_56
timestamp 1626908933
transform 1 0 11232 0 -1 18648
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1017
timestamp 1626908933
transform 1 0 11376 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_229
timestamp 1626908933
transform 1 0 11376 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_949
timestamp 1626908933
transform 1 0 11376 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_181
timestamp 1626908933
transform 1 0 11376 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1013
timestamp 1626908933
transform 1 0 11664 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_225
timestamp 1626908933
transform 1 0 11664 0 1 18167
box -29 -23 29 23
use M1M2_PR  M1M2_PR_944
timestamp 1626908933
transform 1 0 11664 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_176
timestamp 1626908933
transform 1 0 11664 0 1 18167
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_76
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_346
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_76
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_346
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_76
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_346
timestamp 1626908933
transform 1 0 12600 0 1 17982
box -200 -49 200 49
use L1M1_PR  L1M1_PR_642
timestamp 1626908933
transform 1 0 12432 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1430
timestamp 1626908933
transform 1 0 12432 0 1 18389
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_2
timestamp 1626908933
transform 1 0 11328 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_12
timestamp 1626908933
transform 1 0 11328 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_12
timestamp 1626908933
transform 1 0 11328 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_2
timestamp 1626908933
transform 1 0 11328 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_34
timestamp 1626908933
transform 1 0 12480 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_293
timestamp 1626908933
transform 1 0 12480 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_390
timestamp 1626908933
transform 1 0 12768 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_959
timestamp 1626908933
transform 1 0 12768 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_37
timestamp 1626908933
transform 1 0 12576 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_405
timestamp 1626908933
transform 1 0 12576 0 -1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_185
timestamp 1626908933
transform 1 0 13104 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_953
timestamp 1626908933
transform 1 0 13104 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_221
timestamp 1626908933
transform 1 0 13296 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_235
timestamp 1626908933
transform 1 0 13200 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1009
timestamp 1626908933
transform 1 0 13296 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1023
timestamp 1626908933
transform 1 0 13200 0 1 18315
box -29 -23 29 23
use M1M2_PR  M1M2_PR_174
timestamp 1626908933
transform 1 0 13488 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_942
timestamp 1626908933
transform 1 0 13488 0 1 18167
box -32 -32 32 32
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_3
timestamp 1626908933
transform 1 0 13152 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_13
timestamp 1626908933
transform 1 0 13152 0 -1 18648
box -38 -49 1190 715
use L1M1_PR  L1M1_PR_1434
timestamp 1626908933
transform 1 0 14352 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_646
timestamp 1626908933
transform 1 0 14352 0 1 18093
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_225
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_513
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_481
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_211
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_481
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_211
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_481
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_211
timestamp 1626908933
transform 1 0 14600 0 1 18648
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_36
timestamp 1626908933
transform 1 0 15072 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_404
timestamp 1626908933
transform 1 0 15072 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_26
timestamp 1626908933
transform 1 0 14976 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_285
timestamp 1626908933
transform 1 0 14976 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_31
timestamp 1626908933
transform 1 0 15072 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_399
timestamp 1626908933
transform 1 0 15072 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_1
timestamp 1626908933
transform 1 0 14304 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  sky130_fd_sc_hs__fill_8_3
timestamp 1626908933
transform 1 0 14304 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_13
timestamp 1626908933
transform 1 0 13152 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_3
timestamp 1626908933
transform 1 0 13152 0 1 18648
box -38 -49 1862 715
use osc_core_VIA7  osc_core_VIA7_331
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_61
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_331
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_61
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_331
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_61
timestamp 1626908933
transform 1 0 16600 0 1 17982
box -200 -49 200 49
use M1M2_PR  M1M2_PR_1359
timestamp 1626908933
transform 1 0 15504 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_591
timestamp 1626908933
transform 1 0 15504 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1051
timestamp 1626908933
transform 1 0 16368 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_263
timestamp 1626908933
transform 1 0 16368 0 1 18167
box -29 -23 29 23
use M1M2_PR  M1M2_PR_215
timestamp 1626908933
transform 1 0 16272 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_983
timestamp 1626908933
transform 1 0 16272 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_266
timestamp 1626908933
transform 1 0 16272 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1054
timestamp 1626908933
transform 1 0 16272 0 1 18315
box -29 -23 29 23
use M2M3_PR  M2M3_PR_33
timestamp 1626908933
transform 1 0 16080 0 1 18337
box -33 -37 33 37
use M2M3_PR  M2M3_PR_92
timestamp 1626908933
transform 1 0 16080 0 1 18337
box -33 -37 33 37
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_382
timestamp 1626908933
transform 1 0 15264 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_952
timestamp 1626908933
transform 1 0 15264 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_6
timestamp 1626908933
transform 1 0 16032 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_16
timestamp 1626908933
transform 1 0 16032 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_381
timestamp 1626908933
transform 1 0 15264 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_951
timestamp 1626908933
transform 1 0 15264 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_358
timestamp 1626908933
transform 1 0 17184 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_726
timestamp 1626908933
transform 1 0 17184 0 -1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_211
timestamp 1626908933
transform 1 0 16656 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_615
timestamp 1626908933
transform 1 0 17232 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_979
timestamp 1626908933
transform 1 0 16656 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1383
timestamp 1626908933
transform 1 0 17232 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_658
timestamp 1626908933
transform 1 0 17232 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1446
timestamp 1626908933
transform 1 0 17232 0 1 18093
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1228
timestamp 1626908933
transform 1 0 17376 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_598
timestamp 1626908933
transform 1 0 17376 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_292
timestamp 1626908933
transform 1 0 17472 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_33
timestamp 1626908933
transform 1 0 17472 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_727
timestamp 1626908933
transform 1 0 17568 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_359
timestamp 1626908933
transform 1 0 17568 0 -1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_975
timestamp 1626908933
transform 1 0 17616 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_207
timestamp 1626908933
transform 1 0 17616 0 1 18167
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1229
timestamp 1626908933
transform 1 0 17760 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_599
timestamp 1626908933
transform 1 0 17760 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_989
timestamp 1626908933
transform 1 0 17808 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_221
timestamp 1626908933
transform 1 0 17808 0 1 18315
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1061
timestamp 1626908933
transform 1 0 17904 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_273
timestamp 1626908933
transform 1 0 17904 0 1 18315
box -29 -23 29 23
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_7
timestamp 1626908933
transform 1 0 17856 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_17
timestamp 1626908933
transform 1 0 17856 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_17
timestamp 1626908933
transform 1 0 17856 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_7
timestamp 1626908933
transform 1 0 17856 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_16
timestamp 1626908933
transform 1 0 16032 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_6
timestamp 1626908933
transform 1 0 16032 0 1 18648
box -38 -49 1862 715
use L1M1_PR  L1M1_PR_1046
timestamp 1626908933
transform 1 0 18000 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_258
timestamp 1626908933
transform 1 0 18000 0 1 18167
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_497
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_209
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_466
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_196
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_466
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_196
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_466
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_196
timestamp 1626908933
transform 1 0 18600 0 1 18648
box -200 -49 200 49
use M1M2_PR  M1M2_PR_584
timestamp 1626908933
transform 1 0 19344 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1352
timestamp 1626908933
transform 1 0 19344 0 1 18093
box -32 -32 32 32
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_0
timestamp 1626908933
transform 1 0 19008 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_9
timestamp 1626908933
transform 1 0 19008 0 -1 18648
box -38 -49 422 715
use M1M2_PR  M1M2_PR_623
timestamp 1626908933
transform 1 0 19056 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1391
timestamp 1626908933
transform 1 0 19056 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_662
timestamp 1626908933
transform 1 0 19056 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1450
timestamp 1626908933
transform 1 0 19056 0 1 18093
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_362
timestamp 1626908933
transform 1 0 19680 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_730
timestamp 1626908933
transform 1 0 19680 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_604
timestamp 1626908933
transform 1 0 19872 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1234
timestamp 1626908933
transform 1 0 19872 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_25
timestamp 1626908933
transform 1 0 19968 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_284
timestamp 1626908933
transform 1 0 19968 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_605
timestamp 1626908933
transform 1 0 20064 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1235
timestamp 1626908933
transform 1 0 20064 0 1 18648
box -38 -49 134 715
use osc_core_VIA7  osc_core_VIA7_316
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_46
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_316
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_46
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_316
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_46
timestamp 1626908933
transform 1 0 20600 0 1 17982
box -200 -49 200 49
use M1M2_PR  M1M2_PR_968
timestamp 1626908933
transform 1 0 20304 0 1 18093
box -32 -32 32 32
use M1M2_PR  M1M2_PR_200
timestamp 1626908933
transform 1 0 20304 0 1 18093
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1038
timestamp 1626908933
transform 1 0 20112 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_250
timestamp 1626908933
transform 1 0 20112 0 1 18093
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1032
timestamp 1626908933
transform 1 0 20496 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_244
timestamp 1626908933
transform 1 0 20496 0 1 18167
box -29 -23 29 23
use M1M2_PR  M1M2_PR_963
timestamp 1626908933
transform 1 0 20496 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_195
timestamp 1626908933
transform 1 0 20496 0 1 18167
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_310
timestamp 1626908933
transform 1 0 19392 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_880
timestamp 1626908933
transform 1 0 19392 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_4
timestamp 1626908933
transform 1 0 20160 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_14
timestamp 1626908933
transform 1 0 20160 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_14
timestamp 1626908933
transform 1 0 20160 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_4
timestamp 1626908933
transform 1 0 20160 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_35
timestamp 1626908933
transform 1 0 21312 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_403
timestamp 1626908933
transform 1 0 21312 0 -1 18648
box -38 -49 230 715
use M1M2_PR  M1M2_PR_191
timestamp 1626908933
transform 1 0 20880 0 1 18167
box -32 -32 32 32
use M1M2_PR  M1M2_PR_959
timestamp 1626908933
transform 1 0 20880 0 1 18167
box -32 -32 32 32
use L1M1_PR  L1M1_PR_650
timestamp 1626908933
transform 1 0 21264 0 1 18389
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1438
timestamp 1626908933
transform 1 0 21264 0 1 18389
box -29 -23 29 23
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_32
timestamp 1626908933
transform 1 0 21888 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_291
timestamp 1626908933
transform 1 0 21888 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_203
timestamp 1626908933
transform 1 0 21936 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_971
timestamp 1626908933
transform 1 0 21936 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_601
timestamp 1626908933
transform 1 0 21840 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1369
timestamp 1626908933
transform 1 0 21840 0 1 18537
box -32 -32 32 32
use L1M1_PR  L1M1_PR_239
timestamp 1626908933
transform 1 0 22128 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_254
timestamp 1626908933
transform 1 0 22032 0 1 18315
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1027
timestamp 1626908933
transform 1 0 22128 0 1 18167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1042
timestamp 1626908933
transform 1 0 22032 0 1 18315
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_813
timestamp 1626908933
transform 1 0 21504 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_244
timestamp 1626908933
transform 1 0 21504 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_5
timestamp 1626908933
transform 1 0 21984 0 -1 18648
box -38 -49 1190 715
use sky130_fd_sc_hs__einvp_4  sky130_fd_sc_hs__einvp_4_15
timestamp 1626908933
transform 1 0 21984 0 -1 18648
box -38 -49 1190 715
use osc_core_VIA5  osc_core_VIA5_181
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_451
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_181
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_451
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_181
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_451
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_193
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_481
timestamp 1626908933
transform 1 0 22600 0 1 18648
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_34
timestamp 1626908933
transform 1 0 23136 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_402
timestamp 1626908933
transform 1 0 23136 0 -1 18648
box -38 -49 230 715
use L1M1_PR  L1M1_PR_654
timestamp 1626908933
transform 1 0 23184 0 1 18241
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1442
timestamp 1626908933
transform 1 0 23184 0 1 18241
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_242
timestamp 1626908933
transform 1 0 23328 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_812
timestamp 1626908933
transform 1 0 23328 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_15
timestamp 1626908933
transform 1 0 21984 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__einvp_8  sky130_fd_sc_hs__einvp_8_5
timestamp 1626908933
transform 1 0 21984 0 1 18648
box -38 -49 1862 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_674
timestamp 1626908933
transform 1 0 23808 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_44
timestamp 1626908933
transform 1 0 23808 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_794
timestamp 1626908933
transform 1 0 23904 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_224
timestamp 1626908933
transform 1 0 23904 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_779
timestamp 1626908933
transform 1 0 24096 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_210
timestamp 1626908933
transform 1 0 24096 0 -1 18648
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_301
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_31
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_301
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_31
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_301
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_31
timestamp 1626908933
transform 1 0 24600 0 1 17982
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_398
timestamp 1626908933
transform 1 0 24672 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_30
timestamp 1626908933
transform 1 0 24672 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_685
timestamp 1626908933
transform 1 0 24480 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_55
timestamp 1626908933
transform 1 0 24480 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_43
timestamp 1626908933
transform 1 0 24864 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_673
timestamp 1626908933
transform 1 0 24864 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_24
timestamp 1626908933
transform 1 0 24960 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_283
timestamp 1626908933
transform 1 0 24960 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_29
timestamp 1626908933
transform 1 0 25056 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_397
timestamp 1626908933
transform 1 0 25056 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_221
timestamp 1626908933
transform 1 0 24576 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_791
timestamp 1626908933
transform 1 0 24576 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_54
timestamp 1626908933
transform 1 0 25344 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_684
timestamp 1626908933
transform 1 0 25344 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_598
timestamp 1626908933
transform 1 0 25968 0 1 18315
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1366
timestamp 1626908933
transform 1 0 25968 0 1 18315
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_199
timestamp 1626908933
transform 1 0 25824 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_769
timestamp 1626908933
transform 1 0 25824 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_195
timestamp 1626908933
transform 1 0 25440 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_764
timestamp 1626908933
transform 1 0 25440 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_175
timestamp 1626908933
transform 1 0 26016 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_744
timestamp 1626908933
transform 1 0 26016 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_202
timestamp 1626908933
transform 1 0 25248 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_772
timestamp 1626908933
transform 1 0 25248 0 1 18648
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_465
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_177
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_436
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_166
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_436
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_166
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_436
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_166
timestamp 1626908933
transform 1 0 26600 0 1 18648
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_672
timestamp 1626908933
transform 1 0 26400 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_42
timestamp 1626908933
transform 1 0 26400 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_683
timestamp 1626908933
transform 1 0 26592 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_53
timestamp 1626908933
transform 1 0 26592 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_599
timestamp 1626908933
transform 1 0 26928 0 1 18537
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1367
timestamp 1626908933
transform 1 0 26928 0 1 18537
box -32 -32 32 32
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_177
timestamp 1626908933
transform 1 0 26688 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_747
timestamp 1626908933
transform 1 0 26688 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_180
timestamp 1626908933
transform 1 0 26496 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_750
timestamp 1626908933
transform 1 0 26496 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_33
timestamp 1626908933
transform 1 0 27552 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_401
timestamp 1626908933
transform 1 0 27552 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_31
timestamp 1626908933
transform 1 0 27456 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_290
timestamp 1626908933
transform 1 0 27456 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_28
timestamp 1626908933
transform 1 0 27264 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_396
timestamp 1626908933
transform 1 0 27264 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_52
timestamp 1626908933
transform 1 0 27744 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_682
timestamp 1626908933
transform 1 0 27744 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_156
timestamp 1626908933
transform 1 0 27840 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_726
timestamp 1626908933
transform 1 0 27840 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_161
timestamp 1626908933
transform 1 0 27456 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_730
timestamp 1626908933
transform 1 0 27456 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_155
timestamp 1626908933
transform 1 0 27840 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_725
timestamp 1626908933
transform 1 0 27840 0 1 18648
box -38 -49 806 715
use osc_core_VIA5  osc_core_VIA5_16
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_286
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_16
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_286
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_16
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_286
timestamp 1626908933
transform 1 0 28600 0 1 17982
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_138
timestamp 1626908933
transform 1 0 28608 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_707
timestamp 1626908933
transform 1 0 28608 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_137
timestamp 1626908933
transform 1 0 28608 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_706
timestamp 1626908933
transform 1 0 28608 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_671
timestamp 1626908933
transform 1 0 28992 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_41
timestamp 1626908933
transform 1 0 28992 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_681
timestamp 1626908933
transform 1 0 28992 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_51
timestamp 1626908933
transform 1 0 28992 0 -1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_604
timestamp 1626908933
transform 1 0 29328 0 1 18241
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1372
timestamp 1626908933
transform 1 0 29328 0 1 18241
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_50
timestamp 1626908933
transform 1 0 29856 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_680
timestamp 1626908933
transform 1 0 29856 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_606
timestamp 1626908933
transform 1 0 29856 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1236
timestamp 1626908933
transform 1 0 29856 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_132
timestamp 1626908933
transform 1 0 29088 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_702
timestamp 1626908933
transform 1 0 29088 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_131
timestamp 1626908933
transform 1 0 29088 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_701
timestamp 1626908933
transform 1 0 29088 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_40
timestamp 1626908933
transform 1 0 30240 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_670
timestamp 1626908933
transform 1 0 30240 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_23
timestamp 1626908933
transform 1 0 29952 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_282
timestamp 1626908933
transform 1 0 29952 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_27
timestamp 1626908933
transform 1 0 30048 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_395
timestamp 1626908933
transform 1 0 30048 0 1 18648
box -38 -49 230 715
use osc_core_VIA5  osc_core_VIA5_151
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_421
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_151
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_421
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_151
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_421
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_161
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_449
timestamp 1626908933
transform 1 0 30600 0 1 18648
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_107
timestamp 1626908933
transform 1 0 30336 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_677
timestamp 1626908933
transform 1 0 30336 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_118
timestamp 1626908933
transform 1 0 29952 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_687
timestamp 1626908933
transform 1 0 29952 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_106
timestamp 1626908933
transform 1 0 30336 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_676
timestamp 1626908933
transform 1 0 30336 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_394
timestamp 1626908933
transform 1 0 31104 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_26
timestamp 1626908933
transform 1 0 31104 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_654
timestamp 1626908933
transform 1 0 31296 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_85
timestamp 1626908933
transform 1 0 31296 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_400
timestamp 1626908933
transform 1 0 31104 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_32
timestamp 1626908933
transform 1 0 31104 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_655
timestamp 1626908933
transform 1 0 31296 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_86
timestamp 1626908933
transform 1 0 31296 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_646
timestamp 1626908933
transform 1 0 31680 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_76
timestamp 1626908933
transform 1 0 31680 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_647
timestamp 1626908933
transform 1 0 31680 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_77
timestamp 1626908933
transform 1 0 31680 0 -1 18648
box -38 -49 806 715
use osc_core_VIA7  osc_core_VIA7_271
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_1
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_271
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_1
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_271
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_1
timestamp 1626908933
transform 1 0 32600 0 1 17982
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_669
timestamp 1626908933
transform 1 0 32448 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_39
timestamp 1626908933
transform 1 0 32448 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_289
timestamp 1626908933
transform 1 0 32448 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_30
timestamp 1626908933
transform 1 0 32448 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_53
timestamp 1626908933
transform 1 0 32544 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_622
timestamp 1626908933
transform 1 0 32544 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_52
timestamp 1626908933
transform 1 0 32544 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_621
timestamp 1626908933
transform 1 0 32544 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_616
timestamp 1626908933
transform 1 0 32928 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_46
timestamp 1626908933
transform 1 0 32928 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_617
timestamp 1626908933
transform 1 0 32928 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_47
timestamp 1626908933
transform 1 0 32928 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_49
timestamp 1626908933
transform 1 0 33696 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_679
timestamp 1626908933
transform 1 0 33696 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_38
timestamp 1626908933
transform 1 0 33696 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_668
timestamp 1626908933
transform 1 0 33696 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_17
timestamp 1626908933
transform 1 0 34176 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_587
timestamp 1626908933
transform 1 0 34176 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_20
timestamp 1626908933
transform 1 0 33792 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_589
timestamp 1626908933
transform 1 0 33792 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_16
timestamp 1626908933
transform 1 0 34176 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_586
timestamp 1626908933
transform 1 0 34176 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_19
timestamp 1626908933
transform 1 0 33792 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_588
timestamp 1626908933
transform 1 0 33792 0 1 18648
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_406
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_136
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_406
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_136
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_406
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_136
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_145
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_433
timestamp 1626908933
transform 1 0 34600 0 1 18648
box -200 -142 200 178
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_731
timestamp 1626908933
transform 1 0 35424 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_363
timestamp 1626908933
transform 1 0 35424 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_570
timestamp 1626908933
transform 1 0 35040 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1
timestamp 1626908933
transform 1 0 35040 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_281
timestamp 1626908933
transform 1 0 34944 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_22
timestamp 1626908933
transform 1 0 34944 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_571
timestamp 1626908933
transform 1 0 34944 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1
timestamp 1626908933
transform 1 0 34944 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1237
timestamp 1626908933
transform 1 0 35616 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_607
timestamp 1626908933
transform 1 0 35616 0 1 18648
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1399
timestamp 1626908933
transform 1 0 48 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_631
timestamp 1626908933
transform 1 0 48 0 1 19425
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_667
timestamp 1626908933
transform 1 0 288 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_37
timestamp 1626908933
transform 1 0 288 0 -1 19980
box -38 -49 134 715
use M2M3_PR  M2M3_PR_99
timestamp 1626908933
transform 1 0 48 0 1 18825
box -33 -37 33 37
use M2M3_PR  M2M3_PR_40
timestamp 1626908933
transform 1 0 48 0 1 18825
box -33 -37 33 37
use M1M2_PR  M1M2_PR_163
timestamp 1626908933
transform 1 0 1104 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_931
timestamp 1626908933
transform 1 0 1104 0 1 18907
box -32 -32 32 32
use osc_core_VIA5  osc_core_VIA5_120
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_390
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_120
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_390
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_120
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_390
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_417
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_129
timestamp 1626908933
transform 1 0 600 0 1 19314
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_566
timestamp 1626908933
transform 1 0 768 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1136
timestamp 1626908933
transform 1 0 768 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_563
timestamp 1626908933
transform 1 0 384 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1132
timestamp 1626908933
transform 1 0 384 0 -1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_997
timestamp 1626908933
transform 1 0 1200 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_993
timestamp 1626908933
transform 1 0 1200 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_209
timestamp 1626908933
transform 1 0 1200 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_205
timestamp 1626908933
transform 1 0 1200 0 1 19055
box -29 -23 29 23
use M1M2_PR  M1M2_PR_926
timestamp 1626908933
transform 1 0 1296 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_158
timestamp 1626908933
transform 1 0 1296 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_393
timestamp 1626908933
transform 1 0 1536 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_25
timestamp 1626908933
transform 1 0 1536 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1122
timestamp 1626908933
transform 1 0 1728 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_552
timestamp 1626908933
transform 1 0 1728 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_537
timestamp 1626908933
transform 1 0 2688 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1106
timestamp 1626908933
transform 1 0 2688 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_36
timestamp 1626908933
transform 1 0 2592 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_666
timestamp 1626908933
transform 1 0 2592 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_21
timestamp 1626908933
transform 1 0 2496 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_280
timestamp 1626908933
transform 1 0 2496 0 -1 19980
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1423
timestamp 1626908933
transform 1 0 2832 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_635
timestamp 1626908933
transform 1 0 2832 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_936
timestamp 1626908933
transform 1 0 2928 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_168
timestamp 1626908933
transform 1 0 2928 0 1 18907
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1002
timestamp 1626908933
transform 1 0 3024 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_214
timestamp 1626908933
transform 1 0 3024 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_989
timestamp 1626908933
transform 1 0 3024 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_201
timestamp 1626908933
transform 1 0 3024 0 1 19055
box -29 -23 29 23
use M1M2_PR  M1M2_PR_925
timestamp 1626908933
transform 1 0 3216 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_157
timestamp 1626908933
transform 1 0 3216 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_0
timestamp 1626908933
transform 1 0 3072 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_5
timestamp 1626908933
transform 1 0 3072 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_140
timestamp 1626908933
transform -1 0 4992 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_60
timestamp 1626908933
transform -1 0 4992 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_732
timestamp 1626908933
transform 1 0 3936 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_364
timestamp 1626908933
transform 1 0 3936 0 -1 19980
box -38 -49 230 715
use M2M3_PR  M2M3_PR_98
timestamp 1626908933
transform 1 0 4560 0 1 18825
box -33 -37 33 37
use M2M3_PR  M2M3_PR_39
timestamp 1626908933
transform 1 0 4560 0 1 18825
box -33 -37 33 37
use osc_core_VIA7  osc_core_VIA7_375
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_105
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_375
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_105
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_375
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_105
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_401
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_113
timestamp 1626908933
transform 1 0 4600 0 1 19314
box -200 -142 200 178
use L1M1_PR  L1M1_PR_639
timestamp 1626908933
transform 1 0 4656 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1427
timestamp 1626908933
transform 1 0 4656 0 1 18907
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_24
timestamp 1626908933
transform 1 0 4992 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_392
timestamp 1626908933
transform 1 0 4992 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_35
timestamp 1626908933
transform 1 0 5184 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_665
timestamp 1626908933
transform 1 0 5184 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_231
timestamp 1626908933
transform 1 0 5808 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_999
timestamp 1626908933
transform 1 0 5808 0 1 18759
box -32 -32 32 32
use L1M1_PR  L1M1_PR_287
timestamp 1626908933
transform 1 0 5712 0 1 18759
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1075
timestamp 1626908933
transform 1 0 5712 0 1 18759
box -29 -23 29 23
use M1M2_PR  M1M2_PR_226
timestamp 1626908933
transform 1 0 6000 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_994
timestamp 1626908933
transform 1 0 6000 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_497
timestamp 1626908933
transform 1 0 6048 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1066
timestamp 1626908933
transform 1 0 6048 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_519
timestamp 1626908933
transform 1 0 5280 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1089
timestamp 1626908933
transform 1 0 5280 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_124
timestamp 1626908933
transform 1 0 6432 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_44
timestamp 1626908933
transform 1 0 6432 0 -1 19980
box -38 -49 902 715
use M1M2_PR  M1M2_PR_1397
timestamp 1626908933
transform 1 0 6192 0 1 19425
box -32 -32 32 32
use M1M2_PR  M1M2_PR_629
timestamp 1626908933
transform 1 0 6192 0 1 19425
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1069
timestamp 1626908933
transform 1 0 6096 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_281
timestamp 1626908933
transform 1 0 6096 0 1 19055
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_365
timestamp 1626908933
transform 1 0 7296 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_733
timestamp 1626908933
transform 1 0 7296 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_279
timestamp 1626908933
transform 1 0 7488 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_20
timestamp 1626908933
transform 1 0 7488 0 -1 19980
box -38 -49 134 715
use L1M1_PR  L1M1_PR_1455
timestamp 1626908933
transform 1 0 7536 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_667
timestamp 1626908933
transform 1 0 7536 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1401
timestamp 1626908933
transform 1 0 7440 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_633
timestamp 1626908933
transform 1 0 7440 0 1 18907
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1078
timestamp 1626908933
transform 1 0 7728 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_290
timestamp 1626908933
transform 1 0 7728 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1003
timestamp 1626908933
transform 1 0 7632 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_235
timestamp 1626908933
transform 1 0 7632 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1407
timestamp 1626908933
transform 1 0 7824 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_993
timestamp 1626908933
transform 1 0 7824 0 1 19055
box -32 -32 32 32
use M1M2_PR  M1M2_PR_639
timestamp 1626908933
transform 1 0 7824 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_225
timestamp 1626908933
transform 1 0 7824 0 1 19055
box -32 -32 32 32
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_4
timestamp 1626908933
transform 1 0 7584 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_9
timestamp 1626908933
transform 1 0 7584 0 -1 19980
box -38 -49 902 715
use L1M1_PR  L1M1_PR_276
timestamp 1626908933
transform 1 0 7920 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1064
timestamp 1626908933
transform 1 0 7920 0 1 19055
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_385
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_97
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_360
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_90
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_360
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_90
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_360
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_90
timestamp 1626908933
transform 1 0 8600 0 1 19314
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_664
timestamp 1626908933
transform 1 0 8448 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_34
timestamp 1626908933
transform 1 0 8448 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_487
timestamp 1626908933
transform 1 0 8544 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1057
timestamp 1626908933
transform 1 0 8544 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_663
timestamp 1626908933
transform 1 0 9312 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_33
timestamp 1626908933
transform 1 0 9312 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1030
timestamp 1626908933
transform 1 0 9408 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_461
timestamp 1626908933
transform 1 0 9408 0 -1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1459
timestamp 1626908933
transform 1 0 9360 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_671
timestamp 1626908933
transform 1 0 9360 0 1 18907
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1044
timestamp 1626908933
transform 1 0 9792 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_474
timestamp 1626908933
transform 1 0 9792 0 -1 19980
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1344
timestamp 1626908933
transform 1 0 10320 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_576
timestamp 1626908933
transform 1 0 10320 0 1 18759
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_32
timestamp 1626908933
transform 1 0 10560 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_662
timestamp 1626908933
transform 1 0 10560 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_180
timestamp 1626908933
transform 1 0 11376 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_948
timestamp 1626908933
transform 1 0 11376 0 1 18759
box -32 -32 32 32
use L1M1_PR  L1M1_PR_231
timestamp 1626908933
transform 1 0 11280 0 1 18759
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1019
timestamp 1626908933
transform 1 0 11280 0 1 18759
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_453
timestamp 1626908933
transform 1 0 11040 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_1023
timestamp 1626908933
transform 1 0 11040 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_438
timestamp 1626908933
transform 1 0 10656 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1007
timestamp 1626908933
transform 1 0 10656 0 -1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_175
timestamp 1626908933
transform 1 0 11664 0 1 18833
box -32 -32 32 32
use M1M2_PR  M1M2_PR_943
timestamp 1626908933
transform 1 0 11664 0 1 18833
box -32 -32 32 32
use L1M1_PR  L1M1_PR_224
timestamp 1626908933
transform 1 0 11664 0 1 18833
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1012
timestamp 1626908933
transform 1 0 11664 0 1 18833
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_23
timestamp 1626908933
transform 1 0 11808 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_391
timestamp 1626908933
transform 1 0 11808 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_31
timestamp 1626908933
transform 1 0 12000 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_661
timestamp 1626908933
transform 1 0 12000 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_413
timestamp 1626908933
transform 1 0 12096 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_982
timestamp 1626908933
transform 1 0 12096 0 -1 19980
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_369
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_81
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_345
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_75
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_345
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_75
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_345
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_75
timestamp 1626908933
transform 1 0 12600 0 1 19314
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_19
timestamp 1626908933
transform 1 0 12480 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_278
timestamp 1626908933
transform 1 0 12480 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_389
timestamp 1626908933
transform 1 0 12768 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_958
timestamp 1626908933
transform 1 0 12768 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_22
timestamp 1626908933
transform 1 0 12576 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_390
timestamp 1626908933
transform 1 0 12576 0 -1 19980
box -38 -49 230 715
use M1M2_PR  M1M2_PR_184
timestamp 1626908933
transform 1 0 13104 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_952
timestamp 1626908933
transform 1 0 13104 0 1 18759
box -32 -32 32 32
use L1M1_PR  L1M1_PR_233
timestamp 1626908933
transform 1 0 13296 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_643
timestamp 1626908933
transform 1 0 13104 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1021
timestamp 1626908933
transform 1 0 13296 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1431
timestamp 1626908933
transform 1 0 13104 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_569
timestamp 1626908933
transform 1 0 13296 0 1 19129
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1337
timestamp 1626908933
transform 1 0 13296 0 1 19129
box -32 -32 32 32
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_1
timestamp 1626908933
transform 1 0 13152 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_6
timestamp 1626908933
transform 1 0 13152 0 -1 19980
box -38 -49 902 715
use M1M2_PR  M1M2_PR_173
timestamp 1626908933
transform 1 0 13488 0 1 19129
box -32 -32 32 32
use M1M2_PR  M1M2_PR_941
timestamp 1626908933
transform 1 0 13488 0 1 19129
box -32 -32 32 32
use L1M1_PR  L1M1_PR_220
timestamp 1626908933
transform 1 0 13488 0 1 19129
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1008
timestamp 1626908933
transform 1 0 13488 0 1 19129
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_21
timestamp 1626908933
transform 1 0 14016 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_389
timestamp 1626908933
transform 1 0 14016 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_30
timestamp 1626908933
transform 1 0 14208 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_660
timestamp 1626908933
transform 1 0 14208 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_409
timestamp 1626908933
transform 1 0 14304 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_979
timestamp 1626908933
transform 1 0 14304 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_659
timestamp 1626908933
transform 1 0 15072 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_29
timestamp 1626908933
transform 1 0 15072 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_916
timestamp 1626908933
transform 1 0 15168 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_347
timestamp 1626908933
transform 1 0 15168 0 -1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1435
timestamp 1626908933
transform 1 0 14928 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_647
timestamp 1626908933
transform 1 0 14928 0 1 18907
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_950
timestamp 1626908933
transform 1 0 15552 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_380
timestamp 1626908933
transform 1 0 15552 0 -1 19980
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1057
timestamp 1626908933
transform 1 0 15984 0 1 18833
box -29 -23 29 23
use L1M1_PR  L1M1_PR_269
timestamp 1626908933
transform 1 0 15984 0 1 18833
box -29 -23 29 23
use M1M2_PR  M1M2_PR_982
timestamp 1626908933
transform 1 0 16272 0 1 18833
box -32 -32 32 32
use M1M2_PR  M1M2_PR_214
timestamp 1626908933
transform 1 0 16272 0 1 18833
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_353
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_65
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_330
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_60
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_330
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_60
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_330
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_60
timestamp 1626908933
transform 1 0 16600 0 1 19314
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_388
timestamp 1626908933
transform 1 0 16320 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_20
timestamp 1626908933
transform 1 0 16320 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_658
timestamp 1626908933
transform 1 0 16512 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_28
timestamp 1626908933
transform 1 0 16512 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_210
timestamp 1626908933
transform 1 0 16656 0 1 18981
box -32 -32 32 32
use M1M2_PR  M1M2_PR_978
timestamp 1626908933
transform 1 0 16656 0 1 18981
box -32 -32 32 32
use L1M1_PR  L1M1_PR_261
timestamp 1626908933
transform 1 0 16848 0 1 18981
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1049
timestamp 1626908933
transform 1 0 16848 0 1 18981
box -29 -23 29 23
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_355
timestamp 1626908933
transform 1 0 16608 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_925
timestamp 1626908933
transform 1 0 16608 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_277
timestamp 1626908933
transform 1 0 17376 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_18
timestamp 1626908933
transform 1 0 17376 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_8
timestamp 1626908933
transform 1 0 17472 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_3
timestamp 1626908933
transform 1 0 17472 0 -1 19980
box -38 -49 902 715
use L1M1_PR  L1M1_PR_1447
timestamp 1626908933
transform 1 0 17808 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_659
timestamp 1626908933
transform 1 0 17808 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_987
timestamp 1626908933
transform 1 0 17904 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_219
timestamp 1626908933
transform 1 0 17904 0 1 18907
box -32 -32 32 32
use L1M1_PR  L1M1_PR_257
timestamp 1626908933
transform 1 0 18000 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_271
timestamp 1626908933
transform 1 0 18000 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1045
timestamp 1626908933
transform 1 0 18000 0 1 19055
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1059
timestamp 1626908933
transform 1 0 18000 0 1 18907
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_27
timestamp 1626908933
transform 1 0 18336 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_657
timestamp 1626908933
transform 1 0 18336 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_332
timestamp 1626908933
transform 1 0 18816 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_902
timestamp 1626908933
transform 1 0 18816 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_293
timestamp 1626908933
transform 1 0 18432 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_862
timestamp 1626908933
transform 1 0 18432 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_845
timestamp 1626908933
transform 1 0 19584 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_276
timestamp 1626908933
transform 1 0 19584 0 -1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1451
timestamp 1626908933
transform 1 0 19632 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_663
timestamp 1626908933
transform 1 0 19632 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1394
timestamp 1626908933
transform 1 0 19632 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_626
timestamp 1626908933
transform 1 0 19632 0 1 18907
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_26
timestamp 1626908933
transform 1 0 19968 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_656
timestamp 1626908933
transform 1 0 19968 0 -1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_585
timestamp 1626908933
transform 1 0 20112 0 1 19129
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1353
timestamp 1626908933
transform 1 0 20112 0 1 19129
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1035
timestamp 1626908933
transform 1 0 20304 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_247
timestamp 1626908933
transform 1 0 20304 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_967
timestamp 1626908933
transform 1 0 20304 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_199
timestamp 1626908933
transform 1 0 20304 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_194
timestamp 1626908933
transform 1 0 20496 0 1 19129
box -32 -32 32 32
use M1M2_PR  M1M2_PR_962
timestamp 1626908933
transform 1 0 20496 0 1 19129
box -32 -32 32 32
use L1M1_PR  L1M1_PR_243
timestamp 1626908933
transform 1 0 20496 0 1 19129
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1031
timestamp 1626908933
transform 1 0 20496 0 1 19129
box -29 -23 29 23
use osc_core_VIA5  osc_core_VIA5_45
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_315
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_45
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_315
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_45
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_315
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_49
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_337
timestamp 1626908933
transform 1 0 20600 0 1 19314
box -200 -142 200 178
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_297
timestamp 1626908933
transform 1 0 20064 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_867
timestamp 1626908933
transform 1 0 20064 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_655
timestamp 1626908933
transform 1 0 21024 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_25
timestamp 1626908933
transform 1 0 21024 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_387
timestamp 1626908933
transform 1 0 20832 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_19
timestamp 1626908933
transform 1 0 20832 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_817
timestamp 1626908933
transform 1 0 21120 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_248
timestamp 1626908933
transform 1 0 21120 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_7
timestamp 1626908933
transform 1 0 21504 0 -1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_2
timestamp 1626908933
transform 1 0 21504 0 -1 19980
box -38 -49 902 715
use M1M2_PR  M1M2_PR_600
timestamp 1626908933
transform 1 0 21840 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1368
timestamp 1626908933
transform 1 0 21840 0 1 18907
box -32 -32 32 32
use L1M1_PR  L1M1_PR_651
timestamp 1626908933
transform 1 0 21936 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1439
timestamp 1626908933
transform 1 0 21936 0 1 18907
box -29 -23 29 23
use M1M2_PR  M1M2_PR_202
timestamp 1626908933
transform 1 0 22032 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_970
timestamp 1626908933
transform 1 0 22032 0 1 18907
box -32 -32 32 32
use L1M1_PR  L1M1_PR_252
timestamp 1626908933
transform 1 0 22128 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1040
timestamp 1626908933
transform 1 0 22128 0 1 18907
box -29 -23 29 23
use L1M1_PR  L1M1_PR_238
timestamp 1626908933
transform 1 0 22128 0 1 19129
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1026
timestamp 1626908933
transform 1 0 22128 0 1 19129
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_608
timestamp 1626908933
transform 1 0 22368 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1238
timestamp 1626908933
transform 1 0 22368 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_17
timestamp 1626908933
transform 1 0 22464 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_276
timestamp 1626908933
transform 1 0 22464 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_24
timestamp 1626908933
transform 1 0 22560 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_654
timestamp 1626908933
transform 1 0 22560 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_815
timestamp 1626908933
transform 1 0 22656 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_245
timestamp 1626908933
transform 1 0 22656 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_781
timestamp 1626908933
transform 1 0 23424 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_212
timestamp 1626908933
transform 1 0 23424 0 -1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1361
timestamp 1626908933
transform 1 0 23472 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_593
timestamp 1626908933
transform 1 0 23472 0 1 18759
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_653
timestamp 1626908933
transform 1 0 23808 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_23
timestamp 1626908933
transform 1 0 23808 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_793
timestamp 1626908933
transform 1 0 23904 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_223
timestamp 1626908933
transform 1 0 23904 0 -1 19980
box -38 -49 806 715
use L1M1_PR  L1M1_PR_1443
timestamp 1626908933
transform 1 0 23856 0 1 18833
box -29 -23 29 23
use L1M1_PR  L1M1_PR_655
timestamp 1626908933
transform 1 0 23856 0 1 18833
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_321
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_33
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_300
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_30
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_300
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_30
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_300
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_30
timestamp 1626908933
transform 1 0 24600 0 1 19314
box -200 -49 200 49
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_386
timestamp 1626908933
transform 1 0 24672 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_18
timestamp 1626908933
transform 1 0 24672 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_198
timestamp 1626908933
transform 1 0 24864 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_767
timestamp 1626908933
transform 1 0 24864 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_771
timestamp 1626908933
transform 1 0 25248 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_201
timestamp 1626908933
transform 1 0 25248 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_743
timestamp 1626908933
transform 1 0 26016 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_174
timestamp 1626908933
transform 1 0 26016 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_652
timestamp 1626908933
transform 1 0 26400 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_22
timestamp 1626908933
transform 1 0 26400 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_749
timestamp 1626908933
transform 1 0 26496 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_179
timestamp 1626908933
transform 1 0 26496 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_17
timestamp 1626908933
transform 1 0 27552 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_385
timestamp 1626908933
transform 1 0 27552 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_16
timestamp 1626908933
transform 1 0 27456 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_275
timestamp 1626908933
transform 1 0 27456 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_21
timestamp 1626908933
transform 1 0 27264 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_609
timestamp 1626908933
transform 1 0 27360 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_651
timestamp 1626908933
transform 1 0 27264 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1239
timestamp 1626908933
transform 1 0 27360 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_20
timestamp 1626908933
transform 1 0 27744 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_650
timestamp 1626908933
transform 1 0 27744 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_154
timestamp 1626908933
transform 1 0 27840 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_724
timestamp 1626908933
transform 1 0 27840 0 -1 19980
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_305
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_17
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_15
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_285
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_15
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_285
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_15
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_285
timestamp 1626908933
transform 1 0 28600 0 1 19314
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_136
timestamp 1626908933
transform 1 0 28608 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_705
timestamp 1626908933
transform 1 0 28608 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_649
timestamp 1626908933
transform 1 0 28992 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_19
timestamp 1626908933
transform 1 0 28992 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_700
timestamp 1626908933
transform 1 0 29088 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_130
timestamp 1626908933
transform 1 0 29088 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_648
timestamp 1626908933
transform 1 0 29856 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_18
timestamp 1626908933
transform 1 0 29856 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_686
timestamp 1626908933
transform 1 0 29952 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_117
timestamp 1626908933
transform 1 0 29952 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_675
timestamp 1626908933
transform 1 0 30336 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_105
timestamp 1626908933
transform 1 0 30336 0 -1 19980
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1373
timestamp 1626908933
transform 1 0 30192 0 1 18759
box -32 -32 32 32
use M1M2_PR  M1M2_PR_605
timestamp 1626908933
transform 1 0 30192 0 1 18759
box -32 -32 32 32
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_384
timestamp 1626908933
transform 1 0 31104 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_16
timestamp 1626908933
transform 1 0 31104 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_653
timestamp 1626908933
transform 1 0 31296 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_84
timestamp 1626908933
transform 1 0 31296 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_645
timestamp 1626908933
transform 1 0 31680 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_75
timestamp 1626908933
transform 1 0 31680 0 -1 19980
box -38 -49 806 715
use osc_core_VIA4  osc_core_VIA4_289
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_1
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -142 200 178
use osc_core_VIA7  osc_core_VIA7_270
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_0
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_270
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_0
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_270
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_0
timestamp 1626908933
transform 1 0 32600 0 1 19314
box -200 -49 200 49
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_274
timestamp 1626908933
transform 1 0 32448 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_15
timestamp 1626908933
transform 1 0 32448 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_51
timestamp 1626908933
transform 1 0 32544 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_620
timestamp 1626908933
transform 1 0 32544 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_615
timestamp 1626908933
transform 1 0 32928 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_45
timestamp 1626908933
transform 1 0 32928 0 -1 19980
box -38 -49 806 715
use M1M2_PR  M1M2_PR_1385
timestamp 1626908933
transform 1 0 33456 0 1 18907
box -32 -32 32 32
use M1M2_PR  M1M2_PR_617
timestamp 1626908933
transform 1 0 33456 0 1 18907
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_647
timestamp 1626908933
transform 1 0 33696 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_17
timestamp 1626908933
transform 1 0 33696 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_587
timestamp 1626908933
transform 1 0 33792 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_18
timestamp 1626908933
transform 1 0 33792 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_585
timestamp 1626908933
transform 1 0 34176 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_15
timestamp 1626908933
transform 1 0 34176 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_0
timestamp 1626908933
transform 1 0 34944 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_570
timestamp 1626908933
transform 1 0 34944 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_646
timestamp 1626908933
transform 1 0 384 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_16
timestamp 1626908933
transform 1 0 384 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1131
timestamp 1626908933
transform 1 0 480 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_562
timestamp 1626908933
transform 1 0 480 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_273
timestamp 1626908933
transform 1 0 288 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_14
timestamp 1626908933
transform 1 0 288 0 1 19980
box -38 -49 134 715
use M2M3_PR  M2M3_PR_97
timestamp 1626908933
transform 1 0 48 0 1 19801
box -33 -37 33 37
use M2M3_PR  M2M3_PR_38
timestamp 1626908933
transform 1 0 48 0 1 19801
box -33 -37 33 37
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1124
timestamp 1626908933
transform 1 0 864 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_555
timestamp 1626908933
transform 1 0 864 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1123
timestamp 1626908933
transform 1 0 1248 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_554
timestamp 1626908933
transform 1 0 1248 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1121
timestamp 1626908933
transform 1 0 1632 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_552
timestamp 1626908933
transform 1 0 1632 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1117
timestamp 1626908933
transform 1 0 2016 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_548
timestamp 1626908933
transform 1 0 2016 0 1 19980
box -38 -49 422 715
use osc_core_VIA7  osc_core_VIA7_525
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_255
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_525
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_255
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_525
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_255
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_560
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_272
timestamp 1626908933
transform 1 0 2600 0 1 19980
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_645
timestamp 1626908933
transform 1 0 2400 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_15
timestamp 1626908933
transform 1 0 2400 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_383
timestamp 1626908933
transform 1 0 2592 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_15
timestamp 1626908933
transform 1 0 2592 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1105
timestamp 1626908933
transform 1 0 2784 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_536
timestamp 1626908933
transform 1 0 2784 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_272
timestamp 1626908933
transform 1 0 2496 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_13
timestamp 1626908933
transform 1 0 2496 0 1 19980
box -38 -49 134 715
use L1M1_PR  L1M1_PR_988
timestamp 1626908933
transform 1 0 3216 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_200
timestamp 1626908933
transform 1 0 3216 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_924
timestamp 1626908933
transform 1 0 3216 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_156
timestamp 1626908933
transform 1 0 3216 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1402
timestamp 1626908933
transform 1 0 3216 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_614
timestamp 1626908933
transform 1 0 3216 0 1 19869
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1307
timestamp 1626908933
transform 1 0 3120 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_539
timestamp 1626908933
transform 1 0 3120 0 1 19869
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1103
timestamp 1626908933
transform 1 0 3168 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_534
timestamp 1626908933
transform 1 0 3168 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1096
timestamp 1626908933
transform 1 0 3552 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_527
timestamp 1626908933
transform 1 0 3552 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_141
timestamp 1626908933
transform -1 0 4896 0 1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_61
timestamp 1626908933
transform -1 0 4896 0 1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1240
timestamp 1626908933
transform 1 0 3936 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_610
timestamp 1626908933
transform 1 0 3936 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_139
timestamp 1626908933
transform 1 0 4272 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_907
timestamp 1626908933
transform 1 0 4272 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_137
timestamp 1626908933
transform 1 0 4464 0 1 19721
box -32 -32 32 32
use M1M2_PR  M1M2_PR_905
timestamp 1626908933
transform 1 0 4464 0 1 19721
box -32 -32 32 32
use L1M1_PR  L1M1_PR_174
timestamp 1626908933
transform 1 0 4464 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_962
timestamp 1626908933
transform 1 0 4464 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_756
timestamp 1626908933
transform 1 0 4752 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1524
timestamp 1626908933
transform 1 0 4752 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_781
timestamp 1626908933
transform 1 0 4752 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1569
timestamp 1626908933
transform 1 0 4752 0 1 19647
box -29 -23 29 23
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_611
timestamp 1626908933
transform 1 0 4896 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1241
timestamp 1626908933
transform 1 0 4896 0 1 19980
box -38 -49 134 715
use M2M3_PR  M2M3_PR_37
timestamp 1626908933
transform 1 0 5040 0 1 19801
box -33 -37 33 37
use M2M3_PR  M2M3_PR_96
timestamp 1626908933
transform 1 0 5040 0 1 19801
box -33 -37 33 37
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_14
timestamp 1626908933
transform 1 0 5088 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_382
timestamp 1626908933
transform 1 0 5088 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_12
timestamp 1626908933
transform 1 0 4992 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_271
timestamp 1626908933
transform 1 0 4992 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1075
timestamp 1626908933
transform 1 0 5760 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_506
timestamp 1626908933
transform 1 0 5760 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_644
timestamp 1626908933
transform 1 0 5280 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_14
timestamp 1626908933
transform 1 0 5280 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1078
timestamp 1626908933
transform 1 0 5376 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_509
timestamp 1626908933
transform 1 0 5376 0 1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1507
timestamp 1626908933
transform 1 0 6288 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_739
timestamp 1626908933
transform 1 0 6288 0 1 19647
box -32 -32 32 32
use osc_core_VIA7  osc_core_VIA7_510
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_240
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_510
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_240
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_510
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_240
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -49 200 49
use osc_core_VIA4  osc_core_VIA4_256
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_544
timestamp 1626908933
transform 1 0 6600 0 1 19980
box -200 -142 200 178
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1242
timestamp 1626908933
transform 1 0 6240 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_643
timestamp 1626908933
transform 1 0 6144 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_612
timestamp 1626908933
transform 1 0 6240 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_13
timestamp 1626908933
transform 1 0 6144 0 1 19980
box -38 -49 134 715
use L1M1_PR  L1M1_PR_765
timestamp 1626908933
transform 1 0 6576 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1553
timestamp 1626908933
transform 1 0 6576 0 1 19647
box -29 -23 29 23
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_45
timestamp 1626908933
transform 1 0 6336 0 1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_125
timestamp 1626908933
transform 1 0 6336 0 1 19980
box -38 -49 902 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1243
timestamp 1626908933
transform 1 0 7392 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_613
timestamp 1626908933
transform 1 0 7392 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_734
timestamp 1626908933
transform 1 0 7200 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_366
timestamp 1626908933
transform 1 0 7200 0 1 19980
box -38 -49 230 715
use L1M1_PR  L1M1_PR_882
timestamp 1626908933
transform 1 0 7056 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_94
timestamp 1626908933
transform 1 0 7056 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_850
timestamp 1626908933
transform 1 0 7056 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_82
timestamp 1626908933
transform 1 0 7056 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_543
timestamp 1626908933
transform 1 0 7536 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1311
timestamp 1626908933
transform 1 0 7536 0 1 19869
box -32 -32 32 32
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_11
timestamp 1626908933
transform 1 0 7488 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_270
timestamp 1626908933
transform 1 0 7488 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_224
timestamp 1626908933
transform 1 0 7824 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_992
timestamp 1626908933
transform 1 0 7824 0 1 19647
box -32 -32 32 32
use L1M1_PR  L1M1_PR_277
timestamp 1626908933
transform 1 0 7824 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1065
timestamp 1626908933
transform 1 0 7824 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_618
timestamp 1626908933
transform 1 0 7728 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1406
timestamp 1626908933
transform 1 0 7728 0 1 19869
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_484
timestamp 1626908933
transform 1 0 7584 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1053
timestamp 1626908933
transform 1 0 7584 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1052
timestamp 1626908933
transform 1 0 7968 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_483
timestamp 1626908933
transform 1 0 7968 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1050
timestamp 1626908933
transform 1 0 8352 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1038
timestamp 1626908933
transform 1 0 8736 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_481
timestamp 1626908933
transform 1 0 8352 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_469
timestamp 1626908933
transform 1 0 8736 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1037
timestamp 1626908933
transform 1 0 9120 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_468
timestamp 1626908933
transform 1 0 9120 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1029
timestamp 1626908933
transform 1 0 9504 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_460
timestamp 1626908933
transform 1 0 9504 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1244
timestamp 1626908933
transform 1 0 9888 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_614
timestamp 1626908933
transform 1 0 9888 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_381
timestamp 1626908933
transform 1 0 10080 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_13
timestamp 1626908933
transform 1 0 10080 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_269
timestamp 1626908933
transform 1 0 9984 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_10
timestamp 1626908933
transform 1 0 9984 0 1 19980
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_240
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_528
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_225
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_495
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_225
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_495
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_225
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_495
timestamp 1626908933
transform 1 0 10600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_441
timestamp 1626908933
transform 1 0 10272 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1010
timestamp 1626908933
transform 1 0 10272 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1006
timestamp 1626908933
transform 1 0 10656 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_1005
timestamp 1626908933
transform 1 0 11040 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_437
timestamp 1626908933
transform 1 0 10656 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_436
timestamp 1626908933
transform 1 0 11040 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_990
timestamp 1626908933
transform 1 0 11424 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_421
timestamp 1626908933
transform 1 0 11424 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_642
timestamp 1626908933
transform 1 0 12000 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_12
timestamp 1626908933
transform 1 0 12000 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_380
timestamp 1626908933
transform 1 0 11808 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_12
timestamp 1626908933
transform 1 0 11808 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_981
timestamp 1626908933
transform 1 0 12096 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_412
timestamp 1626908933
transform 1 0 12096 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_268
timestamp 1626908933
transform 1 0 12480 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_9
timestamp 1626908933
transform 1 0 12480 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_641
timestamp 1626908933
transform 1 0 12768 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_11
timestamp 1626908933
transform 1 0 12768 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_379
timestamp 1626908933
transform 1 0 12576 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_11
timestamp 1626908933
transform 1 0 12576 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_957
timestamp 1626908933
transform 1 0 12864 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_388
timestamp 1626908933
transform 1 0 12864 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1403
timestamp 1626908933
transform 1 0 13296 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_615
timestamp 1626908933
transform 1 0 13296 0 1 19869
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_955
timestamp 1626908933
transform 1 0 13248 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_386
timestamp 1626908933
transform 1 0 13248 0 1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1308
timestamp 1626908933
transform 1 0 13392 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_540
timestamp 1626908933
transform 1 0 13392 0 1 19869
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_954
timestamp 1626908933
transform 1 0 13632 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_385
timestamp 1626908933
transform 1 0 13632 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1007
timestamp 1626908933
transform 1 0 13488 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_219
timestamp 1626908933
transform 1 0 13488 0 1 19647
box -29 -23 29 23
use M1M2_PR  M1M2_PR_940
timestamp 1626908933
transform 1 0 13488 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_172
timestamp 1626908933
transform 1 0 13488 0 1 19647
box -32 -32 32 32
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_940
timestamp 1626908933
transform 1 0 14016 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_371
timestamp 1626908933
transform 1 0 14016 0 1 19980
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_224
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_512
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_210
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_480
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_210
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_480
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_210
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_480
timestamp 1626908933
transform 1 0 14600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_367
timestamp 1626908933
transform 1 0 14400 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_936
timestamp 1626908933
transform 1 0 14400 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_8
timestamp 1626908933
transform 1 0 14976 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_267
timestamp 1626908933
transform 1 0 14976 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_615
timestamp 1626908933
transform 1 0 14880 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1245
timestamp 1626908933
transform 1 0 14880 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_10
timestamp 1626908933
transform 1 0 14784 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_640
timestamp 1626908933
transform 1 0 14784 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_9
timestamp 1626908933
transform 1 0 15072 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_639
timestamp 1626908933
transform 1 0 15072 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_346
timestamp 1626908933
transform 1 0 15168 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_915
timestamp 1626908933
transform 1 0 15168 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_914
timestamp 1626908933
transform 1 0 15552 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_345
timestamp 1626908933
transform 1 0 15552 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_638
timestamp 1626908933
transform 1 0 16128 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_8
timestamp 1626908933
transform 1 0 16128 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_378
timestamp 1626908933
transform 1 0 15936 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_10
timestamp 1626908933
transform 1 0 15936 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_910
timestamp 1626908933
transform 1 0 16224 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_891
timestamp 1626908933
transform 1 0 16608 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_341
timestamp 1626908933
transform 1 0 16224 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_322
timestamp 1626908933
transform 1 0 16608 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_886
timestamp 1626908933
transform 1 0 16992 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_317
timestamp 1626908933
transform 1 0 16992 0 1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_977
timestamp 1626908933
transform 1 0 16848 0 1 19573
box -32 -32 32 32
use M1M2_PR  M1M2_PR_209
timestamp 1626908933
transform 1 0 16848 0 1 19573
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1246
timestamp 1626908933
transform 1 0 17376 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_616
timestamp 1626908933
transform 1 0 17376 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_266
timestamp 1626908933
transform 1 0 17472 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_7
timestamp 1626908933
transform 1 0 17472 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1310
timestamp 1626908933
transform 1 0 17520 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_542
timestamp 1626908933
transform 1 0 17520 0 1 19869
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1405
timestamp 1626908933
transform 1 0 17616 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_617
timestamp 1626908933
transform 1 0 17616 0 1 19869
box -29 -23 29 23
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_377
timestamp 1626908933
transform 1 0 17568 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_9
timestamp 1626908933
transform 1 0 17568 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_868
timestamp 1626908933
transform 1 0 17760 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_299
timestamp 1626908933
transform 1 0 17760 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1048
timestamp 1626908933
transform 1 0 17616 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_260
timestamp 1626908933
transform 1 0 17616 0 1 19647
box -29 -23 29 23
use osc_core_VIA4  osc_core_VIA4_208
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_496
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_195
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_465
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_195
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_465
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_195
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_465
timestamp 1626908933
transform 1 0 18600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_298
timestamp 1626908933
transform 1 0 18144 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_867
timestamp 1626908933
transform 1 0 18144 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_861
timestamp 1626908933
transform 1 0 18528 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_852
timestamp 1626908933
transform 1 0 18912 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_292
timestamp 1626908933
transform 1 0 18528 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_283
timestamp 1626908933
transform 1 0 18912 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_851
timestamp 1626908933
transform 1 0 19296 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_282
timestamp 1626908933
transform 1 0 19296 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_376
timestamp 1626908933
transform 1 0 19680 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_8
timestamp 1626908933
transform 1 0 19680 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_6
timestamp 1626908933
transform 1 0 19968 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_265
timestamp 1626908933
transform 1 0 19968 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_617
timestamp 1626908933
transform 1 0 19872 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1247
timestamp 1626908933
transform 1 0 19872 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_196
timestamp 1626908933
transform 1 0 20304 0 1 19647
box -32 -32 32 32
use M1M2_PR  M1M2_PR_964
timestamp 1626908933
transform 1 0 20304 0 1 19647
box -32 -32 32 32
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_7
timestamp 1626908933
transform 1 0 20256 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_637
timestamp 1626908933
transform 1 0 20256 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_7
timestamp 1626908933
transform 1 0 20064 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_375
timestamp 1626908933
transform 1 0 20064 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_833
timestamp 1626908933
transform 1 0 20352 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_832
timestamp 1626908933
transform 1 0 20736 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_264
timestamp 1626908933
transform 1 0 20352 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_263
timestamp 1626908933
transform 1 0 20736 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_816
timestamp 1626908933
transform 1 0 21120 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_247
timestamp 1626908933
transform 1 0 21120 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1404
timestamp 1626908933
transform 1 0 21648 0 1 19869
box -29 -23 29 23
use L1M1_PR  L1M1_PR_616
timestamp 1626908933
transform 1 0 21648 0 1 19869
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_812
timestamp 1626908933
transform 1 0 21504 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_243
timestamp 1626908933
transform 1 0 21504 0 1 19980
box -38 -49 422 715
use L1M1_PR  L1M1_PR_1029
timestamp 1626908933
transform 1 0 21648 0 1 19647
box -29 -23 29 23
use L1M1_PR  L1M1_PR_241
timestamp 1626908933
transform 1 0 21648 0 1 19647
box -29 -23 29 23
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_811
timestamp 1626908933
transform 1 0 21888 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_242
timestamp 1626908933
transform 1 0 21888 0 1 19980
box -38 -49 422 715
use M1M2_PR  M1M2_PR_1309
timestamp 1626908933
transform 1 0 21744 0 1 19869
box -32 -32 32 32
use M1M2_PR  M1M2_PR_541
timestamp 1626908933
transform 1 0 21744 0 1 19869
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_480
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_192
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_180
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_450
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_180
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_450
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_180
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_450
timestamp 1626908933
transform 1 0 22600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_6
timestamp 1626908933
transform 1 0 22272 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_618
timestamp 1626908933
transform 1 0 22368 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_636
timestamp 1626908933
transform 1 0 22272 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1248
timestamp 1626908933
transform 1 0 22368 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_5
timestamp 1626908933
transform 1 0 22464 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_264
timestamp 1626908933
transform 1 0 22464 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_5
timestamp 1626908933
transform 1 0 22560 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_635
timestamp 1626908933
transform 1 0 22560 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_802
timestamp 1626908933
transform 1 0 22656 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_800
timestamp 1626908933
transform 1 0 23040 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_233
timestamp 1626908933
transform 1 0 22656 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_231
timestamp 1626908933
transform 1 0 23040 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_780
timestamp 1626908933
transform 1 0 23424 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_211
timestamp 1626908933
transform 1 0 23424 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_374
timestamp 1626908933
transform 1 0 23808 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_6
timestamp 1626908933
transform 1 0 23808 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_634
timestamp 1626908933
transform 1 0 24000 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_4
timestamp 1626908933
transform 1 0 24000 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_778
timestamp 1626908933
transform 1 0 24096 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_209
timestamp 1626908933
transform 1 0 24096 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1249
timestamp 1626908933
transform 1 0 24864 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_619
timestamp 1626908933
transform 1 0 24864 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_776
timestamp 1626908933
transform 1 0 24480 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_207
timestamp 1626908933
transform 1 0 24480 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_373
timestamp 1626908933
transform 1 0 25056 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_5
timestamp 1626908933
transform 1 0 25056 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_766
timestamp 1626908933
transform 1 0 25248 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_197
timestamp 1626908933
transform 1 0 25248 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_263
timestamp 1626908933
transform 1 0 24960 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_4
timestamp 1626908933
transform 1 0 24960 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_763
timestamp 1626908933
transform 1 0 25632 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_194
timestamp 1626908933
transform 1 0 25632 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_742
timestamp 1626908933
transform 1 0 26016 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_173
timestamp 1626908933
transform 1 0 26016 0 1 19980
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_176
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_464
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_165
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_435
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_165
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_435
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_165
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_435
timestamp 1626908933
transform 1 0 26600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_172
timestamp 1626908933
transform 1 0 26400 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_741
timestamp 1626908933
transform 1 0 26400 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_372
timestamp 1626908933
transform 1 0 27168 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_4
timestamp 1626908933
transform 1 0 27168 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_740
timestamp 1626908933
transform 1 0 26784 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_171
timestamp 1626908933
transform 1 0 26784 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1250
timestamp 1626908933
transform 1 0 27360 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_620
timestamp 1626908933
transform 1 0 27360 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_729
timestamp 1626908933
transform 1 0 27552 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_160
timestamp 1626908933
transform 1 0 27552 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_262
timestamp 1626908933
transform 1 0 27456 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1626908933
transform 1 0 27456 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_633
timestamp 1626908933
transform 1 0 28128 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_3
timestamp 1626908933
transform 1 0 28128 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_371
timestamp 1626908933
transform 1 0 27936 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_3
timestamp 1626908933
transform 1 0 27936 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_726
timestamp 1626908933
transform 1 0 28224 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_157
timestamp 1626908933
transform 1 0 28224 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_704
timestamp 1626908933
transform 1 0 28608 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_135
timestamp 1626908933
transform 1 0 28608 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_703
timestamp 1626908933
transform 1 0 28992 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_134
timestamp 1626908933
transform 1 0 28992 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_696
timestamp 1626908933
transform 1 0 29376 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_127
timestamp 1626908933
transform 1 0 29376 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1251
timestamp 1626908933
transform 1 0 29856 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_632
timestamp 1626908933
transform 1 0 29760 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_621
timestamp 1626908933
transform 1 0 29856 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_2
timestamp 1626908933
transform 1 0 29760 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_261
timestamp 1626908933
transform 1 0 29952 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1626908933
transform 1 0 29952 0 1 19980
box -38 -49 134 715
use osc_core_VIA4  osc_core_VIA4_160
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_448
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_150
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_420
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_150
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_420
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_150
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_420
timestamp 1626908933
transform 1 0 30600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_116
timestamp 1626908933
transform 1 0 30144 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_685
timestamp 1626908933
transform 1 0 30144 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1
timestamp 1626908933
transform 1 0 30048 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_631
timestamp 1626908933
transform 1 0 30048 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_683
timestamp 1626908933
transform 1 0 30528 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_114
timestamp 1626908933
transform 1 0 30528 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_682
timestamp 1626908933
transform 1 0 30912 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_113
timestamp 1626908933
transform 1 0 30912 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_652
timestamp 1626908933
transform 1 0 31296 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_83
timestamp 1626908933
transform 1 0 31296 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_370
timestamp 1626908933
transform 1 0 31680 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_2
timestamp 1626908933
transform 1 0 31680 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_630
timestamp 1626908933
transform 1 0 31872 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_0
timestamp 1626908933
transform 1 0 31872 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_650
timestamp 1626908933
transform 1 0 31968 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_81
timestamp 1626908933
transform 1 0 31968 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1252
timestamp 1626908933
transform 1 0 32352 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_622
timestamp 1626908933
transform 1 0 32352 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_369
timestamp 1626908933
transform 1 0 32544 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_1
timestamp 1626908933
transform 1 0 32544 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_619
timestamp 1626908933
transform 1 0 32736 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_50
timestamp 1626908933
transform 1 0 32736 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_260
timestamp 1626908933
transform 1 0 32448 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1626908933
transform 1 0 32448 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_618
timestamp 1626908933
transform 1 0 33120 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_49
timestamp 1626908933
transform 1 0 33120 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_617
timestamp 1626908933
transform 1 0 33504 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_48
timestamp 1626908933
transform 1 0 33504 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_586
timestamp 1626908933
transform 1 0 33888 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_17
timestamp 1626908933
transform 1 0 33888 0 1 19980
box -38 -49 422 715
use osc_core_VIA4  osc_core_VIA4_144
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_432
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -142 200 178
use osc_core_VIA5  osc_core_VIA5_135
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -49 200 49
use osc_core_VIA5  osc_core_VIA5_405
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_135
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -49 200 49
use osc_core_VIA6  osc_core_VIA6_405
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_135
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -49 200 49
use osc_core_VIA7  osc_core_VIA7_405
timestamp 1626908933
transform 1 0 34600 0 1 19980
box -200 -49 200 49
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_16
timestamp 1626908933
transform 1 0 34272 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_585
timestamp 1626908933
transform 1 0 34272 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1253
timestamp 1626908933
transform 1 0 34848 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_623
timestamp 1626908933
transform 1 0 34848 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_368
timestamp 1626908933
transform 1 0 34656 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_0
timestamp 1626908933
transform 1 0 34656 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_569
timestamp 1626908933
transform 1 0 35040 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_0
timestamp 1626908933
transform 1 0 35040 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_259
timestamp 1626908933
transform 1 0 34944 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0
timestamp 1626908933
transform 1 0 34944 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_735
timestamp 1626908933
transform 1 0 35424 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_367
timestamp 1626908933
transform 1 0 35424 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1254
timestamp 1626908933
transform 1 0 35616 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_624
timestamp 1626908933
transform 1 0 35616 0 1 19980
box -38 -49 134 715
use M1M2_PR  M1M2_PR_1395
timestamp 1626908933
transform 1 0 48 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_627
timestamp 1626908933
transform 1 0 48 0 1 20239
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_128
timestamp 1626908933
transform 1 0 600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_416
timestamp 1626908933
transform 1 0 600 0 1 20553
box -200 -142 200 178
use osc_core_VIA10  osc_core_VIA10_21
timestamp 1626908933
transform 1 0 600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_7
timestamp 1626908933
transform 1 0 600 0 1 20623
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_21
timestamp 1626908933
transform 1 0 600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_7
timestamp 1626908933
transform 1 0 600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_26
timestamp 1626908933
transform 1 0 600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_8
timestamp 1626908933
transform 1 0 600 0 1 20630
box -200 -33 200 33
use osc_core_VIA4  osc_core_VIA4_112
timestamp 1626908933
transform 1 0 4600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_400
timestamp 1626908933
transform 1 0 4600 0 1 20553
box -200 -142 200 178
use L1M1_PR  L1M1_PR_965
timestamp 1626908933
transform 1 0 4368 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_177
timestamp 1626908933
transform 1 0 4368 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_904
timestamp 1626908933
transform 1 0 4464 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_136
timestamp 1626908933
transform 1 0 4464 0 1 20313
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1568
timestamp 1626908933
transform 1 0 4752 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_780
timestamp 1626908933
transform 1 0 4752 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1523
timestamp 1626908933
transform 1 0 4752 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_755
timestamp 1626908933
transform 1 0 4752 0 1 20313
box -32 -32 32 32
use L1M1_PR  L1M1_PR_1554
timestamp 1626908933
transform 1 0 6480 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_766
timestamp 1626908933
transform 1 0 6480 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_1506
timestamp 1626908933
transform 1 0 6288 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_738
timestamp 1626908933
transform 1 0 6288 0 1 20313
box -32 -32 32 32
use osc_core_VIA18  osc_core_VIA18_1
timestamp 1626908933
transform 1 0 4653 0 1 20623
box -147 -26 147 26
use osc_core_VIA18  osc_core_VIA18_0
timestamp 1626908933
transform 1 0 4653 0 1 20623
box -147 -26 147 26
use osc_core_VIA17  osc_core_VIA17_1
timestamp 1626908933
transform 1 0 4653 0 1 20630
box -147 -33 147 33
use osc_core_VIA17  osc_core_VIA17_0
timestamp 1626908933
transform 1 0 4653 0 1 20630
box -147 -33 147 33
use osc_core_VIA8  osc_core_VIA8_25
timestamp 1626908933
transform 1 0 4600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_7
timestamp 1626908933
transform 1 0 4600 0 1 20630
box -200 -33 200 33
use L1M1_PR  L1M1_PR_881
timestamp 1626908933
transform 1 0 7056 0 1 20313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_93
timestamp 1626908933
transform 1 0 7056 0 1 20313
box -29 -23 29 23
use M1M2_PR  M1M2_PR_849
timestamp 1626908933
transform 1 0 7056 0 1 20313
box -32 -32 32 32
use M1M2_PR  M1M2_PR_81
timestamp 1626908933
transform 1 0 7056 0 1 20313
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_96
timestamp 1626908933
transform 1 0 8600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_384
timestamp 1626908933
transform 1 0 8600 0 1 20553
box -200 -142 200 178
use M1M2_PR  M1M2_PR_843
timestamp 1626908933
transform 1 0 9648 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_75
timestamp 1626908933
transform 1 0 9648 0 1 20387
box -32 -32 32 32
use osc_core_VIA10  osc_core_VIA10_20
timestamp 1626908933
transform 1 0 8600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_6
timestamp 1626908933
transform 1 0 8600 0 1 20623
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_20
timestamp 1626908933
transform 1 0 8600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_6
timestamp 1626908933
transform 1 0 8600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_24
timestamp 1626908933
transform 1 0 8600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_6
timestamp 1626908933
transform 1 0 8600 0 1 20630
box -200 -33 200 33
use M1M2_PR  M1M2_PR_71
timestamp 1626908933
transform 1 0 12144 0 1 20387
box -32 -32 32 32
use M1M2_PR  M1M2_PR_839
timestamp 1626908933
transform 1 0 12144 0 1 20387
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_368
timestamp 1626908933
transform 1 0 12600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_80
timestamp 1626908933
transform 1 0 12600 0 1 20553
box -200 -142 200 178
use osc_core_VIA8  osc_core_VIA8_5
timestamp 1626908933
transform 1 0 12600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_23
timestamp 1626908933
transform 1 0 12600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_5
timestamp 1626908933
transform 1 0 12600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_19
timestamp 1626908933
transform 1 0 12600 0 1 20630
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_5
timestamp 1626908933
transform 1 0 12600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_19
timestamp 1626908933
transform 1 0 12600 0 1 20623
box -200 -26 200 26
use osc_core_VIA8  osc_core_VIA8_4
timestamp 1626908933
transform 1 0 16600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_22
timestamp 1626908933
transform 1 0 16600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_4
timestamp 1626908933
transform 1 0 16600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_18
timestamp 1626908933
transform 1 0 16600 0 1 20630
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_4
timestamp 1626908933
transform 1 0 16600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_18
timestamp 1626908933
transform 1 0 16600 0 1 20623
box -200 -26 200 26
use osc_core_VIA4  osc_core_VIA4_352
timestamp 1626908933
transform 1 0 16600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_64
timestamp 1626908933
transform 1 0 16600 0 1 20553
box -200 -142 200 178
use M1M2_PR  M1M2_PR_1393
timestamp 1626908933
transform 1 0 19632 0 1 20239
box -32 -32 32 32
use M1M2_PR  M1M2_PR_625
timestamp 1626908933
transform 1 0 19632 0 1 20239
box -32 -32 32 32
use osc_core_VIA4  osc_core_VIA4_48
timestamp 1626908933
transform 1 0 20600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_336
timestamp 1626908933
transform 1 0 20600 0 1 20553
box -200 -142 200 178
use osc_core_VIA10  osc_core_VIA10_17
timestamp 1626908933
transform 1 0 20600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_3
timestamp 1626908933
transform 1 0 20600 0 1 20623
box -200 -26 200 26
use osc_core_VIA9  osc_core_VIA9_17
timestamp 1626908933
transform 1 0 20600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_3
timestamp 1626908933
transform 1 0 20600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_21
timestamp 1626908933
transform 1 0 20600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_3
timestamp 1626908933
transform 1 0 20600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_2
timestamp 1626908933
transform 1 0 24600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_20
timestamp 1626908933
transform 1 0 24600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_2
timestamp 1626908933
transform 1 0 24600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_16
timestamp 1626908933
transform 1 0 24600 0 1 20630
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_2
timestamp 1626908933
transform 1 0 24600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_16
timestamp 1626908933
transform 1 0 24600 0 1 20623
box -200 -26 200 26
use osc_core_VIA4  osc_core_VIA4_320
timestamp 1626908933
transform 1 0 24600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_32
timestamp 1626908933
transform 1 0 24600 0 1 20553
box -200 -142 200 178
use osc_core_VIA8  osc_core_VIA8_1
timestamp 1626908933
transform 1 0 28600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_19
timestamp 1626908933
transform 1 0 28600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_1
timestamp 1626908933
transform 1 0 28600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_15
timestamp 1626908933
transform 1 0 28600 0 1 20630
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_1
timestamp 1626908933
transform 1 0 28600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_15
timestamp 1626908933
transform 1 0 28600 0 1 20623
box -200 -26 200 26
use osc_core_VIA4  osc_core_VIA4_304
timestamp 1626908933
transform 1 0 28600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_16
timestamp 1626908933
transform 1 0 28600 0 1 20553
box -200 -142 200 178
use osc_core_VIA8  osc_core_VIA8_0
timestamp 1626908933
transform 1 0 32600 0 1 20630
box -200 -33 200 33
use osc_core_VIA8  osc_core_VIA8_18
timestamp 1626908933
transform 1 0 32600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_0
timestamp 1626908933
transform 1 0 32600 0 1 20630
box -200 -33 200 33
use osc_core_VIA9  osc_core_VIA9_14
timestamp 1626908933
transform 1 0 32600 0 1 20630
box -200 -33 200 33
use osc_core_VIA10  osc_core_VIA10_0
timestamp 1626908933
transform 1 0 32600 0 1 20623
box -200 -26 200 26
use osc_core_VIA10  osc_core_VIA10_14
timestamp 1626908933
transform 1 0 32600 0 1 20623
box -200 -26 200 26
use osc_core_VIA4  osc_core_VIA4_288
timestamp 1626908933
transform 1 0 32600 0 1 20553
box -200 -142 200 178
use osc_core_VIA4  osc_core_VIA4_0
timestamp 1626908933
transform 1 0 32600 0 1 20553
box -200 -142 200 178
<< labels >>
rlabel metal2 s 0 23 97 51 4 glob_en
port 1 nsew
rlabel metal2 s 0 467 97 495 4 delay_con_lsb[4]
port 2 nsew
rlabel metal2 s 0 911 97 939 4 delay_con_lsb[3]
port 3 nsew
rlabel metal2 s 0 1429 97 1457 4 delay_con_lsb[2]
port 4 nsew
rlabel metal2 s 0 1873 97 1901 4 delay_con_lsb[1]
port 5 nsew
rlabel metal2 s 0 2391 97 2419 4 delay_con_lsb[0]
port 6 nsew
rlabel metal2 s 0 2835 97 2863 4 delay_con_msb[7]
port 7 nsew
rlabel metal2 s 0 3353 97 3381 4 delay_con_msb[6]
port 8 nsew
rlabel metal2 s 0 3797 97 3825 4 delay_con_msb[5]
port 9 nsew
rlabel metal2 s 0 4315 97 4343 4 delay_con_msb[4]
port 10 nsew
rlabel metal2 s 0 4759 97 4787 4 delay_con_msb[3]
port 11 nsew
rlabel metal2 s 0 5277 97 5305 4 delay_con_msb[2]
port 12 nsew
rlabel metal2 s 0 5721 97 5749 4 delay_con_msb[1]
port 13 nsew
rlabel metal2 s 0 6239 97 6267 4 delay_con_msb[0]
port 14 nsew
rlabel metal2 s 0 6683 97 6711 4 con_perb_1[3]
port 15 nsew
rlabel metal2 s 0 7127 97 7155 4 con_perb_1[2]
port 16 nsew
rlabel metal2 s 0 7645 97 7673 4 con_perb_1[1]
port 17 nsew
rlabel metal2 s 0 8089 97 8117 4 con_perb_1[0]
port 18 nsew
rlabel metal2 s 0 8607 97 8635 4 con_perb_2[3]
port 19 nsew
rlabel metal2 s 0 9051 97 9079 4 con_perb_2[2]
port 20 nsew
rlabel metal2 s 0 9569 97 9597 4 con_perb_2[1]
port 21 nsew
rlabel metal2 s 0 10531 97 10559 4 con_perb_2[0]
port 22 nsew
rlabel metal2 s 0 10975 97 11003 4 con_perb_3[3]
port 23 nsew
rlabel metal2 s 0 11493 97 11521 4 con_perb_3[2]
port 24 nsew
rlabel metal2 s 0 11937 97 11965 4 con_perb_3[1]
port 25 nsew
rlabel metal2 s 0 12455 97 12483 4 con_perb_3[0]
port 26 nsew
rlabel metal2 s 0 12899 97 12927 4 con_perb_4[3]
port 27 nsew
rlabel metal2 s 0 13417 97 13445 4 con_perb_4[2]
port 28 nsew
rlabel metal2 s 0 13861 97 13889 4 con_perb_4[1]
port 29 nsew
rlabel metal2 s 0 14305 97 14333 4 con_perb_4[0]
port 30 nsew
rlabel metal2 s 0 14823 97 14851 4 con_perb_5[3]
port 31 nsew
rlabel metal2 s 0 15267 97 15295 4 con_perb_5[2]
port 32 nsew
rlabel metal2 s 0 15785 97 15813 4 con_perb_5[1]
port 33 nsew
rlabel metal2 s 0 16229 97 16257 4 con_perb_5[0]
port 34 nsew
rlabel metal2 s 0 10013 97 10041 4 ref_clk
port 35 nsew
rlabel metal2 s 0 16747 97 16775 4 pi1_l[3]
port 36 nsew
rlabel metal2 s 0 17191 97 17219 4 pi1_l[2]
port 37 nsew
rlabel metal2 s 0 17709 97 17737 4 pi1_l[1]
port 38 nsew
rlabel metal2 s 0 18153 97 18181 4 pi1_l[0]
port 39 nsew
rlabel metal2 s 0 18671 97 18699 4 pi1_r[3]
port 40 nsew
rlabel metal2 s 0 19115 97 19143 4 pi1_r[2]
port 41 nsew
rlabel metal2 s 0 19633 97 19661 4 pi1_r[1]
port 42 nsew
rlabel metal2 s 0 20077 97 20105 4 pi1_r[0]
port 43 nsew
rlabel metal2 s 0 20595 97 20623 4 pi2_l[3]
port 44 nsew
rlabel metal2 s 35938 0 35966 97 4 pi2_l[2]
port 45 nsew
rlabel metal2 s 35170 0 35198 97 4 pi2_l[1]
port 46 nsew
rlabel metal2 s 34306 0 34334 97 4 pi2_l[0]
port 47 nsew
rlabel metal2 s 33442 0 33470 97 4 pi2_r[3]
port 48 nsew
rlabel metal2 s 32674 0 32702 97 4 pi2_r[2]
port 49 nsew
rlabel metal2 s 31810 0 31838 97 4 pi2_r[1]
port 50 nsew
rlabel metal2 s 30946 0 30974 97 4 pi2_r[0]
port 51 nsew
rlabel metal2 s 30178 0 30206 97 4 pi3_l[3]
port 52 nsew
rlabel metal2 s 29314 0 29342 97 4 pi3_l[2]
port 53 nsew
rlabel metal2 s 28450 0 28478 97 4 pi3_l[1]
port 54 nsew
rlabel metal2 s 27682 0 27710 97 4 pi3_l[0]
port 55 nsew
rlabel metal2 s 26818 0 26846 97 4 pi3_r[3]
port 56 nsew
rlabel metal2 s 25954 0 25982 97 4 pi3_r[2]
port 57 nsew
rlabel metal2 s 25090 0 25118 97 4 pi3_r[1]
port 58 nsew
rlabel metal2 s 24322 0 24350 97 4 pi3_r[0]
port 59 nsew
rlabel metal2 s 23458 0 23486 97 4 pi4_l[3]
port 60 nsew
rlabel metal2 s 22594 0 22622 97 4 pi4_l[2]
port 61 nsew
rlabel metal2 s 21826 0 21854 97 4 pi4_l[1]
port 62 nsew
rlabel metal2 s 20962 0 20990 97 4 pi4_l[0]
port 63 nsew
rlabel metal2 s 20098 0 20126 97 4 pi4_r[3]
port 64 nsew
rlabel metal2 s 19330 0 19358 97 4 pi4_r[2]
port 65 nsew
rlabel metal2 s 18466 0 18494 97 4 pi4_r[1]
port 66 nsew
rlabel metal2 s 17602 0 17630 97 4 pi4_r[0]
port 67 nsew
rlabel metal2 s 16738 0 16766 97 4 pi5_l[3]
port 68 nsew
rlabel metal2 s 15970 0 15998 97 4 pi5_l[2]
port 69 nsew
rlabel metal2 s 15106 0 15134 97 4 pi5_l[1]
port 70 nsew
rlabel metal2 s 14242 0 14270 97 4 pi5_l[0]
port 71 nsew
rlabel metal2 s 13474 0 13502 97 4 pi5_r[3]
port 72 nsew
rlabel metal2 s 12610 0 12638 97 4 pi5_r[2]
port 73 nsew
rlabel metal2 s 11746 0 11774 97 4 pi5_r[1]
port 74 nsew
rlabel metal2 s 10978 0 11006 97 4 pi5_r[0]
port 75 nsew
rlabel metal2 s 4450 20549 4478 20646 4 osc_000
port 76 nsew
rlabel metal2 s 8098 20549 8126 20646 4 osc_036
port 77 nsew
rlabel metal2 s 15106 20549 15134 20646 4 osc_072
port 78 nsew
rlabel metal2 s 19330 20549 19358 20646 4 osc_108
port 79 nsew
rlabel metal2 s 12130 20549 12158 20646 4 osc_144
port 80 nsew
rlabel metal2 s 5890 0 5918 97 4 inj_en
port 81 nsew
rlabel metal2 s 18082 0 18110 97 4 inj_out
port 82 nsew
rlabel metal2 s 18178 0 18206 97 4 osc_hold
port 83 nsew
rlabel metal2 s 7522 20549 7550 20646 4 p1
port 84 nsew
rlabel metal2 s 17506 20549 17534 20646 4 p2
port 85 nsew
rlabel metal2 s 21730 20549 21758 20646 4 p3
port 86 nsew
rlabel metal2 s 13378 20549 13406 20646 4 p4
port 87 nsew
rlabel metal2 s 3106 20549 3134 20646 4 p5
port 88 nsew
rlabel metal1 s 0 -49 98 49 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 -49 36000 49 4 DVSS:
port 89 nsew
rlabel metal1 s 0 1283 98 1381 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 1283 36000 1381 4 DVSS:
port 89 nsew
rlabel metal1 s 0 2615 98 2713 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 2615 36000 2713 4 DVSS:
port 89 nsew
rlabel metal1 s 0 3947 98 4045 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 3947 36000 4045 4 DVSS:
port 89 nsew
rlabel metal1 s 0 5279 98 5377 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 5279 36000 5377 4 DVSS:
port 89 nsew
rlabel metal1 s 0 6611 98 6709 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 6611 36000 6709 4 DVSS:
port 89 nsew
rlabel metal1 s 0 7943 98 8041 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 7943 36000 8041 4 DVSS:
port 89 nsew
rlabel metal1 s 0 9275 98 9373 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 9275 36000 9373 4 DVSS:
port 89 nsew
rlabel metal1 s 0 10607 98 10705 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 10607 36000 10705 4 DVSS:
port 89 nsew
rlabel metal1 s 0 11939 98 12037 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 11939 36000 12037 4 DVSS:
port 89 nsew
rlabel metal1 s 0 13271 98 13369 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 13271 36000 13369 4 DVSS:
port 89 nsew
rlabel metal1 s 0 14603 98 14701 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 14603 36000 14701 4 DVSS:
port 89 nsew
rlabel metal1 s 0 15935 98 16033 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 15935 36000 16033 4 DVSS:
port 89 nsew
rlabel metal1 s 0 17267 98 17365 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 17267 36000 17365 4 DVSS:
port 89 nsew
rlabel metal1 s 0 18599 98 18697 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 18599 36000 18697 4 DVSS:
port 89 nsew
rlabel metal1 s 0 19931 98 20029 4 DVSS:
port 89 nsew
rlabel metal1 s 35902 19931 36000 20029 4 DVSS:
port 89 nsew
rlabel metal1 s 0 617 98 715 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 617 36000 715 4 DVDD:
port 90 nsew
rlabel metal1 s 0 1949 98 2047 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 1949 36000 2047 4 DVDD:
port 90 nsew
rlabel metal1 s 0 3281 98 3379 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 3281 36000 3379 4 DVDD:
port 90 nsew
rlabel metal1 s 0 4613 98 4711 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 4613 36000 4711 4 DVDD:
port 90 nsew
rlabel metal1 s 0 5945 98 6043 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 5945 36000 6043 4 DVDD:
port 90 nsew
rlabel metal1 s 0 7277 98 7375 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 7277 36000 7375 4 DVDD:
port 90 nsew
rlabel metal1 s 0 8609 98 8707 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 8609 36000 8707 4 DVDD:
port 90 nsew
rlabel metal1 s 0 9941 98 10039 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 9941 36000 10039 4 DVDD:
port 90 nsew
rlabel metal1 s 0 11273 98 11371 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 11273 36000 11371 4 DVDD:
port 90 nsew
rlabel metal1 s 0 12605 98 12703 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 12605 36000 12703 4 DVDD:
port 90 nsew
rlabel metal1 s 0 13937 98 14035 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 13937 36000 14035 4 DVDD:
port 90 nsew
rlabel metal1 s 0 15269 98 15367 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 15269 36000 15367 4 DVDD:
port 90 nsew
rlabel metal1 s 0 16601 98 16699 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 16601 36000 16699 4 DVDD:
port 90 nsew
rlabel metal1 s 0 17933 98 18031 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 17933 36000 18031 4 DVDD:
port 90 nsew
rlabel metal1 s 0 19265 98 19363 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 19265 36000 19363 4 DVDD:
port 90 nsew
rlabel metal1 s 0 20597 98 20695 4 DVDD:
port 90 nsew
rlabel metal1 s 35902 20597 36000 20695 4 DVDD:
port 90 nsew
rlabel metal4 s 3452 6660 3452 6660 4 osc_000
port 76 nsew
rlabel metal4 s 7964 6660 7964 6660 4 osc_036
port 77 nsew
rlabel metal4 s 14012 6660 14012 6660 4 osc_144
port 80 nsew
rlabel metal4 s 17852 6660 17852 6660 4 osc_072
port 78 nsew
rlabel metal4 s 22076 6660 22076 6660 4 osc_108
port 79 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 91 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 92 nsew
rlabel metal2 s 48 37 48 37 4 glob_en
port 1 nsew
rlabel metal2 s 48 481 48 481 4 delay_con_lsb[4]
port 2 nsew
rlabel metal2 s 48 925 48 925 4 delay_con_lsb[3]
port 3 nsew
rlabel metal2 s 48 1443 48 1443 4 delay_con_lsb[2]
port 4 nsew
rlabel metal2 s 48 1887 48 1887 4 delay_con_lsb[1]
port 5 nsew
rlabel metal2 s 48 2405 48 2405 4 delay_con_lsb[0]
port 6 nsew
rlabel metal2 s 48 2849 48 2849 4 delay_con_msb[7]
port 7 nsew
rlabel metal2 s 48 3367 48 3367 4 delay_con_msb[6]
port 8 nsew
rlabel metal2 s 48 3811 48 3811 4 delay_con_msb[5]
port 9 nsew
rlabel metal2 s 48 4329 48 4329 4 delay_con_msb[4]
port 10 nsew
rlabel metal2 s 48 4773 48 4773 4 delay_con_msb[3]
port 11 nsew
rlabel metal2 s 48 5291 48 5291 4 delay_con_msb[2]
port 12 nsew
rlabel metal2 s 48 5735 48 5735 4 delay_con_msb[1]
port 13 nsew
rlabel metal2 s 48 6253 48 6253 4 delay_con_msb[0]
port 14 nsew
rlabel metal2 s 48 6697 48 6697 4 con_perb_1[3]
port 15 nsew
rlabel metal2 s 48 7141 48 7141 4 con_perb_1[2]
port 16 nsew
rlabel metal2 s 48 7659 48 7659 4 con_perb_1[1]
port 17 nsew
rlabel metal2 s 48 8103 48 8103 4 con_perb_1[0]
port 18 nsew
rlabel metal2 s 48 8621 48 8621 4 con_perb_2[3]
port 19 nsew
rlabel metal2 s 48 9065 48 9065 4 con_perb_2[2]
port 20 nsew
rlabel metal2 s 48 9583 48 9583 4 con_perb_2[1]
port 21 nsew
rlabel metal2 s 48 10545 48 10545 4 con_perb_2[0]
port 22 nsew
rlabel metal2 s 48 10989 48 10989 4 con_perb_3[3]
port 23 nsew
rlabel metal2 s 48 11507 48 11507 4 con_perb_3[2]
port 24 nsew
rlabel metal2 s 48 11951 48 11951 4 con_perb_3[1]
port 25 nsew
rlabel metal2 s 48 12469 48 12469 4 con_perb_3[0]
port 26 nsew
rlabel metal2 s 48 12913 48 12913 4 con_perb_4[3]
port 27 nsew
rlabel metal2 s 48 13431 48 13431 4 con_perb_4[2]
port 28 nsew
rlabel metal2 s 48 13875 48 13875 4 con_perb_4[1]
port 29 nsew
rlabel metal2 s 48 14319 48 14319 4 con_perb_4[0]
port 30 nsew
rlabel metal2 s 48 14837 48 14837 4 con_perb_5[3]
port 31 nsew
rlabel metal2 s 48 15281 48 15281 4 con_perb_5[2]
port 32 nsew
rlabel metal2 s 48 15799 48 15799 4 con_perb_5[1]
port 33 nsew
rlabel metal2 s 48 16243 48 16243 4 con_perb_5[0]
port 34 nsew
rlabel metal2 s 48 10027 48 10027 4 ref_clk
port 35 nsew
rlabel metal2 s 48 16761 48 16761 4 pi1_l[3]
port 36 nsew
rlabel metal2 s 48 17205 48 17205 4 pi1_l[2]
port 37 nsew
rlabel metal2 s 48 17723 48 17723 4 pi1_l[1]
port 38 nsew
rlabel metal2 s 48 18167 48 18167 4 pi1_l[0]
port 39 nsew
rlabel metal2 s 48 18685 48 18685 4 pi1_r[3]
port 40 nsew
rlabel metal2 s 48 19129 48 19129 4 pi1_r[2]
port 41 nsew
rlabel metal2 s 48 19647 48 19647 4 pi1_r[1]
port 42 nsew
rlabel metal2 s 48 20091 48 20091 4 pi1_r[0]
port 43 nsew
rlabel metal2 s 48 20609 48 20609 4 pi2_l[3]
port 44 nsew
rlabel metal2 s 35952 48 35952 48 4 pi2_l[2]
port 45 nsew
rlabel metal2 s 35184 48 35184 48 4 pi2_l[1]
port 46 nsew
rlabel metal2 s 34320 48 34320 48 4 pi2_l[0]
port 47 nsew
rlabel metal2 s 33456 48 33456 48 4 pi2_r[3]
port 48 nsew
rlabel metal2 s 32688 48 32688 48 4 pi2_r[2]
port 49 nsew
rlabel metal2 s 31824 48 31824 48 4 pi2_r[1]
port 50 nsew
rlabel metal2 s 30960 48 30960 48 4 pi2_r[0]
port 51 nsew
rlabel metal2 s 30192 48 30192 48 4 pi3_l[3]
port 52 nsew
rlabel metal2 s 29328 48 29328 48 4 pi3_l[2]
port 53 nsew
rlabel metal2 s 28464 48 28464 48 4 pi3_l[1]
port 54 nsew
rlabel metal2 s 27696 48 27696 48 4 pi3_l[0]
port 55 nsew
rlabel metal2 s 26832 48 26832 48 4 pi3_r[3]
port 56 nsew
rlabel metal2 s 25968 48 25968 48 4 pi3_r[2]
port 57 nsew
rlabel metal2 s 25104 48 25104 48 4 pi3_r[1]
port 58 nsew
rlabel metal2 s 24336 48 24336 48 4 pi3_r[0]
port 59 nsew
rlabel metal2 s 23472 48 23472 48 4 pi4_l[3]
port 60 nsew
rlabel metal2 s 22608 48 22608 48 4 pi4_l[2]
port 61 nsew
rlabel metal2 s 21840 48 21840 48 4 pi4_l[1]
port 62 nsew
rlabel metal2 s 20976 48 20976 48 4 pi4_l[0]
port 63 nsew
rlabel metal2 s 20112 48 20112 48 4 pi4_r[3]
port 64 nsew
rlabel metal2 s 19344 48 19344 48 4 pi4_r[2]
port 65 nsew
rlabel metal2 s 18480 48 18480 48 4 pi4_r[1]
port 66 nsew
rlabel metal2 s 17616 48 17616 48 4 pi4_r[0]
port 67 nsew
rlabel metal2 s 16752 48 16752 48 4 pi5_l[3]
port 68 nsew
rlabel metal2 s 15984 48 15984 48 4 pi5_l[2]
port 69 nsew
rlabel metal2 s 15120 48 15120 48 4 pi5_l[1]
port 70 nsew
rlabel metal2 s 14256 48 14256 48 4 pi5_l[0]
port 71 nsew
rlabel metal2 s 13488 48 13488 48 4 pi5_r[3]
port 72 nsew
rlabel metal2 s 12624 48 12624 48 4 pi5_r[2]
port 73 nsew
rlabel metal2 s 11760 48 11760 48 4 pi5_r[1]
port 74 nsew
rlabel metal2 s 10992 48 10992 48 4 pi5_r[0]
port 75 nsew
rlabel metal2 s 4464 20597 4464 20597 4 osc_000
port 76 nsew
rlabel metal2 s 8112 20597 8112 20597 4 osc_036
port 77 nsew
rlabel metal2 s 15120 20597 15120 20597 4 osc_072
port 78 nsew
rlabel metal2 s 19344 20597 19344 20597 4 osc_108
port 79 nsew
rlabel metal2 s 12144 20597 12144 20597 4 osc_144
port 80 nsew
rlabel metal2 s 5904 48 5904 48 4 inj_en
port 81 nsew
rlabel metal2 s 18096 48 18096 48 4 inj_out
port 82 nsew
rlabel metal2 s 18192 48 18192 48 4 osc_hold
port 83 nsew
rlabel metal2 s 7536 20597 7536 20597 4 p1
port 84 nsew
rlabel metal2 s 17520 20597 17520 20597 4 p2
port 85 nsew
rlabel metal2 s 21744 20597 21744 20597 4 p3
port 86 nsew
rlabel metal2 s 13392 20597 13392 20597 4 p4
port 87 nsew
rlabel metal2 s 3120 20597 3120 20597 4 p5
port 88 nsew
rlabel metal1 s 49 0 49 0 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 0 35951 0 4 DVSS:
port 89 nsew
rlabel metal1 s 49 1332 49 1332 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 1332 35951 1332 4 DVSS:
port 89 nsew
rlabel metal1 s 49 2664 49 2664 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 2664 35951 2664 4 DVSS:
port 89 nsew
rlabel metal1 s 49 3996 49 3996 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 3996 35951 3996 4 DVSS:
port 89 nsew
rlabel metal1 s 49 5328 49 5328 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 5328 35951 5328 4 DVSS:
port 89 nsew
rlabel metal1 s 49 6660 49 6660 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 6660 35951 6660 4 DVSS:
port 89 nsew
rlabel metal1 s 49 7992 49 7992 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 7992 35951 7992 4 DVSS:
port 89 nsew
rlabel metal1 s 49 9324 49 9324 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 9324 35951 9324 4 DVSS:
port 89 nsew
rlabel metal1 s 49 10656 49 10656 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 10656 35951 10656 4 DVSS:
port 89 nsew
rlabel metal1 s 49 11988 49 11988 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 11988 35951 11988 4 DVSS:
port 89 nsew
rlabel metal1 s 49 13320 49 13320 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 13320 35951 13320 4 DVSS:
port 89 nsew
rlabel metal1 s 49 14652 49 14652 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 14652 35951 14652 4 DVSS:
port 89 nsew
rlabel metal1 s 49 15984 49 15984 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 15984 35951 15984 4 DVSS:
port 89 nsew
rlabel metal1 s 49 17316 49 17316 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 17316 35951 17316 4 DVSS:
port 89 nsew
rlabel metal1 s 49 18648 49 18648 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 18648 35951 18648 4 DVSS:
port 89 nsew
rlabel metal1 s 49 19980 49 19980 4 DVSS:
port 89 nsew
rlabel metal1 s 35951 19980 35951 19980 4 DVSS:
port 89 nsew
rlabel metal1 s 49 666 49 666 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 666 35951 666 4 DVDD:
port 90 nsew
rlabel metal1 s 49 1998 49 1998 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 1998 35951 1998 4 DVDD:
port 90 nsew
rlabel metal1 s 49 3330 49 3330 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 3330 35951 3330 4 DVDD:
port 90 nsew
rlabel metal1 s 49 4662 49 4662 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 4662 35951 4662 4 DVDD:
port 90 nsew
rlabel metal1 s 49 5994 49 5994 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 5994 35951 5994 4 DVDD:
port 90 nsew
rlabel metal1 s 49 7326 49 7326 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 7326 35951 7326 4 DVDD:
port 90 nsew
rlabel metal1 s 49 8658 49 8658 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 8658 35951 8658 4 DVDD:
port 90 nsew
rlabel metal1 s 49 9990 49 9990 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 9990 35951 9990 4 DVDD:
port 90 nsew
rlabel metal1 s 49 11322 49 11322 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 11322 35951 11322 4 DVDD:
port 90 nsew
rlabel metal1 s 49 12654 49 12654 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 12654 35951 12654 4 DVDD:
port 90 nsew
rlabel metal1 s 49 13986 49 13986 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 13986 35951 13986 4 DVDD:
port 90 nsew
rlabel metal1 s 49 15318 49 15318 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 15318 35951 15318 4 DVDD:
port 90 nsew
rlabel metal1 s 49 16650 49 16650 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 16650 35951 16650 4 DVDD:
port 90 nsew
rlabel metal1 s 49 17982 49 17982 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 17982 35951 17982 4 DVDD:
port 90 nsew
rlabel metal1 s 49 19314 49 19314 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 19314 35951 19314 4 DVDD:
port 90 nsew
rlabel metal1 s 49 20646 49 20646 4 DVDD:
port 90 nsew
rlabel metal1 s 35951 20646 35951 20646 4 DVDD:
port 90 nsew
rlabel metal4 s 3452 6660 3452 6660 4 osc_000
port 76 nsew
rlabel metal4 s 7964 6660 7964 6660 4 osc_036
port 77 nsew
rlabel metal4 s 14012 6660 14012 6660 4 osc_144
port 80 nsew
rlabel metal4 s 17852 6660 17852 6660 4 osc_072
port 78 nsew
rlabel metal4 s 22076 6660 22076 6660 4 osc_108
port 79 nsew
rlabel metal1 s 0 -49 0 -49 4 DVSS
port 91 nsew
rlabel metal1 s 0 617 0 617 4 DVDD
port 92 nsew
<< properties >>
string path 560.400 327.275 560.400 330.225 
<< end >>
