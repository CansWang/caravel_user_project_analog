magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< metal2 >>
rect -147 28 147 33
rect -147 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 147 28
rect -147 -33 147 -28
<< via2 >>
rect -108 -28 -52 28
rect -28 -28 28 28
rect 52 -28 108 28
<< metal3 >>
rect -147 28 147 33
rect -147 -28 -108 28
rect -52 -28 -28 28
rect 28 -28 52 28
rect 108 -28 147 28
rect -147 -33 147 -28
<< end >>
