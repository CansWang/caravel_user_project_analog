magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 0 0 672 49
<< scpmos >>
rect 85 464 115 592
rect 286 368 316 592
rect 376 368 406 592
rect 466 368 496 592
rect 556 368 586 592
<< nmoslvt >>
rect 87 74 117 158
rect 288 74 318 222
rect 374 74 404 222
rect 460 74 490 222
rect 547 74 577 222
<< ndiff >>
rect 231 210 288 222
rect 231 176 243 210
rect 277 176 288 210
rect 30 133 87 158
rect 30 99 42 133
rect 76 99 87 133
rect 30 74 87 99
rect 117 133 174 158
rect 117 99 128 133
rect 162 99 174 133
rect 117 74 174 99
rect 231 120 288 176
rect 231 86 243 120
rect 277 86 288 120
rect 231 74 288 86
rect 318 139 374 222
rect 318 105 329 139
rect 363 105 374 139
rect 318 74 374 105
rect 404 210 460 222
rect 404 176 415 210
rect 449 176 460 210
rect 404 120 460 176
rect 404 86 415 120
rect 449 86 460 120
rect 404 74 460 86
rect 490 199 547 222
rect 490 165 501 199
rect 535 165 547 199
rect 490 74 547 165
rect 577 132 627 222
rect 577 120 637 132
rect 577 86 588 120
rect 622 86 637 120
rect 577 74 637 86
<< pdiff >>
rect 27 580 85 592
rect 27 546 38 580
rect 72 546 85 580
rect 27 510 85 546
rect 27 476 38 510
rect 72 476 85 510
rect 27 464 85 476
rect 115 580 173 592
rect 115 546 128 580
rect 162 546 173 580
rect 115 510 173 546
rect 115 476 128 510
rect 162 476 173 510
rect 115 464 173 476
rect 227 580 286 592
rect 227 546 239 580
rect 273 546 286 580
rect 227 497 286 546
rect 227 463 239 497
rect 273 463 286 497
rect 227 414 286 463
rect 227 380 239 414
rect 273 380 286 414
rect 227 368 286 380
rect 316 580 376 592
rect 316 546 329 580
rect 363 546 376 580
rect 316 482 376 546
rect 316 448 329 482
rect 363 448 376 482
rect 316 368 376 448
rect 406 580 466 592
rect 406 546 419 580
rect 453 546 466 580
rect 406 497 466 546
rect 406 463 419 497
rect 453 463 466 497
rect 406 414 466 463
rect 406 380 419 414
rect 453 380 466 414
rect 406 368 466 380
rect 496 547 556 592
rect 496 513 509 547
rect 543 513 556 547
rect 496 479 556 513
rect 496 445 509 479
rect 543 445 556 479
rect 496 411 556 445
rect 496 377 509 411
rect 543 377 556 411
rect 496 368 556 377
rect 586 580 645 592
rect 586 546 599 580
rect 633 546 645 580
rect 586 497 645 546
rect 586 463 599 497
rect 633 463 645 497
rect 586 414 645 463
rect 586 380 599 414
rect 633 380 645 414
rect 586 368 645 380
<< ndiffc >>
rect 243 176 277 210
rect 42 99 76 133
rect 128 99 162 133
rect 243 86 277 120
rect 329 105 363 139
rect 415 176 449 210
rect 415 86 449 120
rect 501 165 535 199
rect 588 86 622 120
<< pdiffc >>
rect 38 546 72 580
rect 38 476 72 510
rect 128 546 162 580
rect 128 476 162 510
rect 239 546 273 580
rect 239 463 273 497
rect 239 380 273 414
rect 329 546 363 580
rect 329 448 363 482
rect 419 546 453 580
rect 419 463 453 497
rect 419 380 453 414
rect 509 513 543 547
rect 509 445 543 479
rect 509 377 543 411
rect 599 546 633 580
rect 599 463 633 497
rect 599 380 633 414
<< poly >>
rect 82 607 409 637
rect 85 592 115 607
rect 286 592 316 607
rect 376 592 406 607
rect 466 592 496 618
rect 556 592 586 618
rect 85 449 115 464
rect 82 426 117 449
rect 44 410 117 426
rect 44 376 60 410
rect 94 376 117 410
rect 44 342 117 376
rect 286 342 316 368
rect 376 342 406 368
rect 466 353 496 368
rect 556 353 586 368
rect 44 308 60 342
rect 94 308 117 342
rect 44 274 117 308
rect 44 240 60 274
rect 94 240 117 274
rect 166 314 232 330
rect 166 280 182 314
rect 216 294 232 314
rect 216 280 404 294
rect 166 264 404 280
rect 463 274 499 353
rect 553 310 589 353
rect 547 294 651 310
rect 547 274 601 294
rect 44 224 117 240
rect 87 158 117 224
rect 288 222 318 264
rect 374 222 404 264
rect 460 260 601 274
rect 635 260 651 294
rect 460 244 651 260
rect 460 222 490 244
rect 547 222 577 244
rect 87 48 117 74
rect 288 48 318 74
rect 374 48 404 74
rect 460 48 490 74
rect 547 48 577 74
<< polycont >>
rect 60 376 94 410
rect 60 308 94 342
rect 60 240 94 274
rect 182 280 216 314
rect 601 260 635 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 22 580 72 649
rect 22 546 38 580
rect 22 510 72 546
rect 22 476 38 510
rect 22 460 72 476
rect 112 580 178 596
rect 112 546 128 580
rect 162 546 178 580
rect 112 510 178 546
rect 112 476 128 510
rect 162 476 178 510
rect 112 460 178 476
rect 25 410 110 426
rect 25 376 60 410
rect 94 376 110 410
rect 25 342 110 376
rect 25 308 60 342
rect 94 308 110 342
rect 25 274 110 308
rect 25 240 60 274
rect 94 240 110 274
rect 25 224 110 240
rect 144 330 178 460
rect 223 580 280 596
rect 223 546 239 580
rect 273 546 280 580
rect 223 497 280 546
rect 223 463 239 497
rect 273 463 280 497
rect 223 414 280 463
rect 316 580 363 649
rect 316 546 329 580
rect 316 482 363 546
rect 316 448 329 482
rect 316 432 363 448
rect 403 581 649 615
rect 403 580 459 581
rect 403 546 419 580
rect 453 546 459 580
rect 593 580 649 581
rect 403 497 459 546
rect 403 463 419 497
rect 453 463 459 497
rect 223 380 239 414
rect 273 398 280 414
rect 403 414 459 463
rect 403 398 419 414
rect 273 380 419 398
rect 453 380 459 414
rect 223 364 459 380
rect 493 513 509 547
rect 543 513 559 547
rect 493 479 559 513
rect 493 445 509 479
rect 543 445 559 479
rect 493 411 559 445
rect 493 377 509 411
rect 543 377 559 411
rect 493 364 559 377
rect 593 546 599 580
rect 633 546 649 580
rect 593 497 649 546
rect 593 463 599 497
rect 633 463 649 497
rect 593 414 649 463
rect 593 380 599 414
rect 633 380 649 414
rect 593 364 649 380
rect 144 314 232 330
rect 144 280 182 314
rect 216 280 232 314
rect 144 264 232 280
rect 144 162 178 264
rect 26 133 76 162
rect 26 99 42 133
rect 26 17 76 99
rect 112 133 178 162
rect 112 99 128 133
rect 162 99 178 133
rect 112 70 178 99
rect 227 210 449 230
rect 493 226 551 364
rect 227 176 243 210
rect 277 196 415 210
rect 227 120 277 176
rect 227 86 243 120
rect 227 70 277 86
rect 313 139 379 158
rect 313 105 329 139
rect 363 105 379 139
rect 313 17 379 105
rect 415 120 449 176
rect 485 199 551 226
rect 485 165 501 199
rect 535 165 551 199
rect 485 154 551 165
rect 585 294 651 310
rect 585 260 601 294
rect 635 260 651 294
rect 585 162 651 260
rect 449 86 588 120
rect 622 86 640 120
rect 415 70 640 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvn_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 TE_B
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 TE_B
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Z
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Z
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Z
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Z
<< properties >>
string FIXED_BBOX 0 0 672 666
<< end >>
