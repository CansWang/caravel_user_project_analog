magic
tech sky130A
magscale 1 2
timestamp 1626908933
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 0 0 864 49
<< scpmos >>
rect 86 368 116 592
rect 178 368 208 592
rect 276 368 306 592
rect 376 368 406 592
rect 468 368 498 592
rect 558 368 588 592
rect 658 368 688 592
rect 748 368 778 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
rect 370 74 400 222
rect 484 74 514 222
rect 647 74 677 222
rect 736 74 766 222
<< ndiff >>
rect 27 162 84 222
rect 27 128 39 162
rect 73 128 84 162
rect 27 74 84 128
rect 114 184 170 222
rect 114 150 125 184
rect 159 150 170 184
rect 114 116 170 150
rect 114 82 125 116
rect 159 82 170 116
rect 114 74 170 82
rect 200 176 270 222
rect 200 142 225 176
rect 259 142 270 176
rect 200 74 270 142
rect 300 116 370 222
rect 300 82 325 116
rect 359 82 370 116
rect 300 74 370 82
rect 400 116 484 222
rect 400 82 425 116
rect 459 82 484 116
rect 400 74 484 82
rect 514 116 647 222
rect 514 82 525 116
rect 559 82 602 116
rect 636 82 647 116
rect 514 74 647 82
rect 677 184 736 222
rect 677 150 691 184
rect 725 150 736 184
rect 677 74 736 150
rect 766 210 837 222
rect 766 176 791 210
rect 825 176 837 210
rect 766 120 837 176
rect 766 86 791 120
rect 825 86 837 120
rect 766 74 837 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 178 592
rect 116 546 129 580
rect 163 546 178 580
rect 116 499 178 546
rect 116 465 129 499
rect 163 465 178 499
rect 116 368 178 465
rect 208 580 276 592
rect 208 546 229 580
rect 263 546 276 580
rect 208 503 276 546
rect 208 469 229 503
rect 263 469 276 503
rect 208 425 276 469
rect 208 391 229 425
rect 263 391 276 425
rect 208 368 276 391
rect 306 580 376 592
rect 306 546 319 580
rect 353 546 376 580
rect 306 508 376 546
rect 306 474 319 508
rect 353 474 376 508
rect 306 368 376 474
rect 406 576 468 592
rect 406 542 420 576
rect 454 542 468 576
rect 406 508 468 542
rect 406 474 420 508
rect 454 474 468 508
rect 406 440 468 474
rect 406 406 420 440
rect 454 406 468 440
rect 406 368 468 406
rect 498 546 558 592
rect 498 512 511 546
rect 545 512 558 546
rect 498 478 558 512
rect 498 444 511 478
rect 545 444 558 478
rect 498 410 558 444
rect 498 376 511 410
rect 545 376 558 410
rect 498 368 558 376
rect 588 584 658 592
rect 588 550 611 584
rect 645 550 658 584
rect 588 514 658 550
rect 588 480 611 514
rect 645 480 658 514
rect 588 446 658 480
rect 588 412 611 446
rect 645 412 658 446
rect 588 368 658 412
rect 688 584 748 592
rect 688 550 701 584
rect 735 550 748 584
rect 688 516 748 550
rect 688 482 701 516
rect 735 482 748 516
rect 688 368 748 482
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 510 837 546
rect 778 476 791 510
rect 825 476 837 510
rect 778 440 837 476
rect 778 406 791 440
rect 825 406 837 440
rect 778 368 837 406
<< ndiffc >>
rect 39 128 73 162
rect 125 150 159 184
rect 125 82 159 116
rect 225 142 259 176
rect 325 82 359 116
rect 425 82 459 116
rect 525 82 559 116
rect 602 82 636 116
rect 691 150 725 184
rect 791 176 825 210
rect 791 86 825 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 465 163 499
rect 229 546 263 580
rect 229 469 263 503
rect 229 391 263 425
rect 319 546 353 580
rect 319 474 353 508
rect 420 542 454 576
rect 420 474 454 508
rect 420 406 454 440
rect 511 512 545 546
rect 511 444 545 478
rect 511 376 545 410
rect 611 550 645 584
rect 611 480 645 514
rect 611 412 645 446
rect 701 550 735 584
rect 701 482 735 516
rect 791 546 825 580
rect 791 476 825 510
rect 791 406 825 440
<< poly >>
rect 86 592 116 618
rect 178 592 208 618
rect 276 592 306 618
rect 376 592 406 618
rect 468 592 498 618
rect 558 592 588 618
rect 658 592 688 618
rect 748 592 778 618
rect 86 353 116 368
rect 178 353 208 368
rect 276 353 306 368
rect 376 353 406 368
rect 468 353 498 368
rect 558 353 588 368
rect 658 353 688 368
rect 748 353 778 368
rect 83 310 119 353
rect 21 294 119 310
rect 175 336 211 353
rect 273 336 309 353
rect 175 320 309 336
rect 175 300 191 320
rect 21 260 37 294
rect 71 260 119 294
rect 21 244 119 260
rect 170 286 191 300
rect 225 286 259 320
rect 293 286 309 320
rect 373 310 409 353
rect 465 310 501 353
rect 555 310 591 353
rect 655 336 691 353
rect 745 336 781 353
rect 655 320 781 336
rect 170 270 309 286
rect 357 294 423 310
rect 84 222 114 244
rect 170 222 200 270
rect 270 222 300 270
rect 357 260 373 294
rect 407 260 423 294
rect 357 244 423 260
rect 465 294 599 310
rect 655 300 731 320
rect 465 260 481 294
rect 515 260 549 294
rect 583 260 599 294
rect 465 244 599 260
rect 647 286 731 300
rect 765 286 781 320
rect 647 270 781 286
rect 370 222 400 244
rect 484 222 514 244
rect 647 222 677 270
rect 736 222 766 270
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
rect 370 48 400 74
rect 484 48 514 74
rect 647 48 677 74
rect 736 48 766 74
<< polycont >>
rect 37 260 71 294
rect 191 286 225 320
rect 259 286 293 320
rect 373 260 407 294
rect 481 260 515 294
rect 549 260 583 294
rect 731 286 765 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 424 73 463
rect 113 580 179 649
rect 113 546 129 580
rect 163 546 179 580
rect 113 499 179 546
rect 113 465 129 499
rect 163 465 179 499
rect 113 458 179 465
rect 213 580 279 596
rect 213 546 229 580
rect 263 546 279 580
rect 213 503 279 546
rect 213 469 229 503
rect 263 469 279 503
rect 213 425 279 469
rect 319 580 369 649
rect 353 546 369 580
rect 319 508 369 546
rect 353 474 369 508
rect 319 458 369 474
rect 403 584 651 615
rect 403 581 611 584
rect 403 576 455 581
rect 403 542 420 576
rect 454 542 455 576
rect 595 550 611 581
rect 645 550 651 584
rect 403 508 455 542
rect 403 474 420 508
rect 454 474 455 508
rect 213 424 229 425
rect 23 414 229 424
rect 23 380 39 414
rect 73 391 229 414
rect 263 424 279 425
rect 403 440 455 474
rect 403 424 420 440
rect 263 406 420 424
rect 454 406 455 440
rect 263 391 455 406
rect 73 390 455 391
rect 495 546 561 547
rect 495 512 511 546
rect 545 512 561 546
rect 495 478 561 512
rect 495 444 511 478
rect 545 444 561 478
rect 495 410 561 444
rect 595 514 651 550
rect 595 480 611 514
rect 645 480 651 514
rect 685 584 751 649
rect 685 550 701 584
rect 735 550 751 584
rect 685 516 751 550
rect 685 482 701 516
rect 735 482 751 516
rect 685 480 751 482
rect 785 580 841 596
rect 785 546 791 580
rect 825 546 841 580
rect 785 510 841 546
rect 595 446 651 480
rect 785 476 791 510
rect 825 476 841 510
rect 785 446 841 476
rect 595 412 611 446
rect 645 440 841 446
rect 645 412 791 440
rect 23 364 73 380
rect 495 376 511 410
rect 545 378 561 410
rect 775 406 791 412
rect 825 406 841 440
rect 775 390 841 406
rect 545 376 667 378
rect 121 320 309 356
rect 495 344 667 376
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 121 286 191 320
rect 225 286 259 320
rect 293 286 309 320
rect 357 294 423 310
rect 21 252 87 260
rect 357 260 373 294
rect 407 260 423 294
rect 357 252 423 260
rect 21 218 423 252
rect 465 294 599 310
rect 465 260 481 294
rect 515 260 549 294
rect 583 260 599 294
rect 465 236 599 260
rect 633 252 667 344
rect 701 320 839 356
rect 701 286 731 320
rect 765 286 839 320
rect 633 218 841 252
rect 775 210 841 218
rect 23 162 73 184
rect 23 128 39 162
rect 23 17 73 128
rect 109 150 125 184
rect 159 150 175 184
rect 109 116 175 150
rect 209 176 691 184
rect 209 142 225 176
rect 259 150 691 176
rect 725 150 741 184
rect 259 142 275 150
rect 209 119 275 142
rect 686 134 741 150
rect 775 176 791 210
rect 825 176 841 210
rect 775 120 841 176
rect 109 82 125 116
rect 159 85 175 116
rect 309 85 325 116
rect 159 82 325 85
rect 359 82 375 116
rect 109 51 375 82
rect 409 82 425 116
rect 459 82 475 116
rect 409 17 475 82
rect 509 82 525 116
rect 559 82 602 116
rect 636 85 652 116
rect 775 86 791 120
rect 825 86 841 120
rect 775 85 841 86
rect 636 82 841 85
rect 509 51 841 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a31oi_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A3
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 Y
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
rlabel comment s 0 0 0 0 4 a31oi_2
flabel pwell s 432 24 432 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 432 641 432 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 432 641 432 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 432 24 432 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A2
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A2
flabel locali s 816 333 816 333 0 FreeSans 340 0 0 0 A1
flabel locali s 48 259 48 259 0 FreeSans 340 0 0 0 A3
flabel locali s 816 111 816 111 0 FreeSans 340 0 0 0 Y
flabel locali s 816 185 816 185 0 FreeSans 340 0 0 0 Y
flabel locali s 528 259 528 259 0 FreeSans 340 0 0 0 B1
rlabel comment s 0 0 0 0 4 a31oi_2
flabel pwell s 432 24 432 24 0 FreeSans 200 0 0 0 VNB
flabel nwell s 432 641 432 641 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 432 641 432 641 0 FreeSans 340 0 0 0 VPWR
flabel metal1 s 432 24 432 24 0 FreeSans 340 0 0 0 VGND
flabel locali s 144 333 144 333 0 FreeSans 340 0 0 0 A2
flabel locali s 240 333 240 333 0 FreeSans 340 0 0 0 A2
flabel locali s 816 333 816 333 0 FreeSans 340 0 0 0 A1
flabel locali s 48 259 48 259 0 FreeSans 340 0 0 0 A3
flabel locali s 816 111 816 111 0 FreeSans 340 0 0 0 Y
flabel locali s 816 185 816 185 0 FreeSans 340 0 0 0 Y
flabel locali s 528 259 528 259 0 FreeSans 340 0 0 0 B1
<< properties >>
string FIXED_BBOX 0 0 864 666
<< end >>
